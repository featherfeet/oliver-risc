`include "gpu_defines.v"

module gpu(
    // Clock and reset signals.
    input CLOCK_50,                           // 50 MHz clock used as a base clock for communications between the CPU and GPU.
    input reset,                              // Reset (active-high).
    // VGA signals.
    input VGA_CLK,                            // 25 (technically should be 25.175) MHz clock for VGA pixels.
    output wire [3:0] VGA_R,                  // VGA red pin (4-bit resistor DAC).
    output wire [3:0] VGA_G,                  // VGA green pin (4-bit resistor DAC).
    output wire [3:0] VGA_B,                  // VGA blue pin (4-bit resistor DAC).
    output wire VGA_HS,                       // VGA h-sync signal.
    output wire VGA_VS,                       // VGA v-sync signal.
    // CPU interface signals.
    input[$clog2(`GPU_TEXT_BUFFER_LENGTH) - 1:0] cell_to_access, // The index of the character cell to read/write.
    input write_enable, // Set high by the CPU to write character_to_write to text_buffer[cell_to_access]. If low, then the character at text_buffer[cell_to_access] is read out into the character_read output.
    input [7:0] character_to_write, // Used by the CPU to write a character to a location in the text buffer.
    output reg [7:0] character_read // Used to send a character read from the text buffer back to the CPU.
);

integer i;

// Buffer holding the text that is being displayed on-screen. Each cell in the array is a byte (8 bits) storing an ASCII character. The first `GPU_TEXT_DISPLAY_COLUMNS cells are the first row of text, the second `GPU_TEXT_DISPLAY_COLUMNS cells are the second row of text, and so on.
reg[7:0] text_buffer[`GPU_TEXT_BUFFER_LENGTH - 1:0];

// Create a VGA controller with 25 MHz pixel clock.
wire blanking;
wire[9:0] pixel_x;
wire[8:0] pixel_y;
vga640x480 vga(.i_clk(CLOCK_50),
               .i_pix_stb(VGA_CLK),
               .i_rst(~reset),
               .o_hs(VGA_HS),
               .o_vs(VGA_VS),
               .o_blanking(blanking),
               .o_x(pixel_x),
               .o_y(pixel_y));

// Registers for tracking the coordinates of the current pixel being drawn within the current character cell.
reg[$clog2(`GPU_CHARACTER_CELL_WIDTH) - 1:0] character_cell_x; // Units: pixels, Range: 0 to character_cell_width - 1
reg[$clog2(`GPU_CHARACTER_CELL_HEIGHT) - 1:0] character_cell_y; // Units: pixels, Range: 0 to character_cell_height - 1
// Register for tracking the current character cell's location in the text buffer.
reg[$clog2(`GPU_TEXT_BUFFER_LENGTH) - 1:0] current_character_cell; // Units: character cells, Range: 0 to `GPU_TEXT_BUFFER_LENGTH - 1
// Register for tracking the current character cell's location on the screen.
reg[$clog2(`GPU_TEXT_DISPLAY_COLUMNS) - 1:0] current_column; // Units: character cells, Range: 0 to `GPU_TEXT_DISPLAY_COLUMNS - 1

// Combinational logic for rendering pixels.
wire[7:0] current_character; // The character currently being drawn.
wire current_pixel_value; // The value (on or off) of the pixel currently being rendered. Generated by the font_rom module.
assign current_character = text_buffer[current_character_cell]; // The current character is selected from the text buffer using the row and column counters.
// If we're in VGA blanking, then switch off the VGA color pins. Otherwise, use current_pixel_value to set the VGA color pins' values.
assign VGA_R = blanking ? 4'b0000 : (current_pixel_value ? 4'b1111 : 4'b0000);
assign VGA_G = blanking ? 4'b0000 : (current_pixel_value ? 4'b1111 : 4'b0000);
assign VGA_B = blanking ? 4'b0000 : (current_pixel_value ? 4'b1111 : 4'b0000);

// Font glyph lookup table, used to render text characters by determining whether the current pixel should be black or white.
font_rom font_glyphs(.character(current_character),
                     .character_cell_x(character_cell_x),
                     .character_cell_y(character_cell_y),
                     .pixel_value(current_pixel_value));

// Sequential logic for letting the CPU access the GPU's text buffer.
always @(posedge CLOCK_50)
begin
    if (reset)
    begin
        for (i = 0; i < `GPU_TEXT_DISPLAY_COLUMNS; i = i + 1)
            text_buffer[i] <= i + 'd33;
        for (i = `GPU_TEXT_DISPLAY_COLUMNS; i < `GPU_TEXT_BUFFER_LENGTH; i = i + 1)
            text_buffer[i] <= 'd0;
    end
    else
    begin
        if (write_enable)
        begin
            $display("Writing character %c to cell %d in GPU text buffer.", character_to_write, cell_to_access);
            text_buffer[cell_to_access] <= character_to_write;
        end
        else
            character_read <= text_buffer[cell_to_access];
    end
end

// Sequential logic for counting pixels, rows, and columns.
always @(posedge VGA_CLK)
begin
    if (reset)
    begin
        character_cell_x <= 'h0;
        character_cell_y <= 'h0;
        current_character_cell <= 'h0;
        current_column <= 'h0;
        $display("In reset.");
    end
    else if (~blanking)
    begin
        if (current_column == `GPU_TEXT_DISPLAY_COLUMNS)
        begin
            character_cell_x <= 'd0;
            current_column <= 'd0;
            if (character_cell_y != `GPU_CHARACTER_CELL_HEIGHT - 'd1)
                current_character_cell <= current_character_cell - `GPU_TEXT_DISPLAY_COLUMNS;
        end
        else
        begin
            if (character_cell_x == `GPU_CHARACTER_CELL_WIDTH - 'd1)
            begin
                character_cell_x <= 'd0;
                current_column <= current_column + 'd1;
                current_character_cell <= current_character_cell + 'd1;
            end
            else
                character_cell_x <= character_cell_x + 'd1;
        end

        if (pixel_x == 0 && pixel_y == 0)
        begin
            character_cell_y <= 'd0;
            current_character_cell <= 'd0;
        end
        else
        begin
            if (character_cell_y == `GPU_CHARACTER_CELL_HEIGHT)
            begin
                character_cell_y <= 'd0;
            end
            else if (pixel_x == `GPU_DISPLAY_WIDTH_PIXELS)
                character_cell_y <= character_cell_y + 'd1;
        end
        //$display("(%d, %d): COL %d, CELL %d", pixel_x, pixel_y, current_column, current_character_cell);
    end
end

endmodule
