// sdram_system.v

// Generated using ACDS version 13.0sp1 232 at 2020.11.22.00:37:50

`timescale 1 ps / 1 ps
module sdram_system (
		output wire [11:0] sdram_controller_addr,  // sdram_controller.addr
		output wire [1:0]  sdram_controller_ba,    //                 .ba
		output wire        sdram_controller_cas_n, //                 .cas_n
		output wire        sdram_controller_cke,   //                 .cke
		output wire        sdram_controller_cs_n,  //                 .cs_n
		inout  wire [15:0] sdram_controller_dq,    //                 .dq
		output wire [1:0]  sdram_controller_dqm,   //                 .dqm
		output wire        sdram_controller_ras_n, //                 .ras_n
		output wire        sdram_controller_we_n,  //                 .we_n
		input  wire        reset_reset_n,          //            reset.reset_n
		input  wire        clk_clk                 //              clk.clk
	);

	wire    rst_controller_reset_out_reset; // rst_controller:reset_out -> new_sdram_controller_0:reset_n

	sdram_system_new_sdram_controller_0 new_sdram_controller_0 (
		.clk            (clk_clk),                         //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset), // reset.reset_n
		.az_addr        (),                                //    s1.address
		.az_be_n        (),                                //      .byteenable_n
		.az_cs          (),                                //      .chipselect
		.az_data        (),                                //      .writedata
		.az_rd_n        (),                                //      .read_n
		.az_wr_n        (),                                //      .write_n
		.za_data        (),                                //      .readdata
		.za_valid       (),                                //      .readdatavalid
		.za_waitrequest (),                                //      .waitrequest
		.zs_addr        (sdram_controller_addr),           //  wire.export
		.zs_ba          (sdram_controller_ba),             //      .export
		.zs_cas_n       (sdram_controller_cas_n),          //      .export
		.zs_cke         (sdram_controller_cke),            //      .export
		.zs_cs_n        (sdram_controller_cs_n),           //      .export
		.zs_dq          (sdram_controller_dq),             //      .export
		.zs_dqm         (sdram_controller_dqm),            //      .export
		.zs_ras_n       (sdram_controller_ras_n),          //      .export
		.zs_we_n        (sdram_controller_we_n)            //      .export
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                 // reset_in0.reset
		.clk        (clk_clk),                        //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req  (),                               // (terminated)
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

endmodule
