// sdram_system.v

// Generated using ACDS version 13.0sp1 232 at 2019.04.04.00:58:52

`timescale 1 ps / 1 ps
module sdram_system (
		input  wire        clk_clk,                   //              clk.clk
		input  wire        reset_reset_n,             //            reset.reset_n
		output wire        vga_clk_clk,               //          vga_clk.clk
		output wire [11:0] sdram_controller_addr,     // sdram_controller.addr
		output wire [1:0]  sdram_controller_ba,       //                 .ba
		output wire        sdram_controller_cas_n,    //                 .cas_n
		output wire        sdram_controller_cke,      //                 .cke
		output wire        sdram_controller_cs_n,     //                 .cs_n
		inout  wire [15:0] sdram_controller_dq,       //                 .dq
		output wire [1:0]  sdram_controller_dqm,      //                 .dqm
		output wire        sdram_controller_ras_n,    //                 .ras_n
		output wire        sdram_controller_we_n,     //                 .we_n
		input  wire [22:0] avalon_bridge_address,     //    avalon_bridge.address
		input  wire [1:0]  avalon_bridge_byte_enable, //                 .byte_enable
		input  wire        avalon_bridge_read,        //                 .read
		input  wire        avalon_bridge_write,       //                 .write
		input  wire [15:0] avalon_bridge_write_data,  //                 .write_data
		output wire        avalon_bridge_acknowledge, //                 .acknowledge
		output wire [15:0] avalon_bridge_read_data    //                 .read_data
	);

	wire         up_clocks_0_sdram_clk_clk;                                                                      // up_clocks_0:SDRAM_CLK -> [crosser:out_clk, crosser_001:in_clk, id_router:clk, new_sdram_controller_0:clk, new_sdram_controller_0_s1_translator:clk, new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:clk, new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, rsp_xbar_demux:clk, rst_controller_001:clk]
	wire         bridge_0_avalon_master_waitrequest;                                                             // bridge_0_avalon_master_translator:av_waitrequest -> bridge_0:avalon_waitrequest
	wire  [22:0] bridge_0_avalon_master_address;                                                                 // bridge_0:avalon_address -> bridge_0_avalon_master_translator:av_address
	wire  [15:0] bridge_0_avalon_master_writedata;                                                               // bridge_0:avalon_writedata -> bridge_0_avalon_master_translator:av_writedata
	wire         bridge_0_avalon_master_write;                                                                   // bridge_0:avalon_write -> bridge_0_avalon_master_translator:av_write
	wire         bridge_0_avalon_master_read;                                                                    // bridge_0:avalon_read -> bridge_0_avalon_master_translator:av_read
	wire  [15:0] bridge_0_avalon_master_readdata;                                                                // bridge_0_avalon_master_translator:av_readdata -> bridge_0:avalon_readdata
	wire   [1:0] bridge_0_avalon_master_byteenable;                                                              // bridge_0:avalon_byteenable -> bridge_0_avalon_master_translator:av_byteenable
	wire         new_sdram_controller_0_s1_translator_avalon_anti_slave_0_waitrequest;                           // new_sdram_controller_0:za_waitrequest -> new_sdram_controller_0_s1_translator:av_waitrequest
	wire  [15:0] new_sdram_controller_0_s1_translator_avalon_anti_slave_0_writedata;                             // new_sdram_controller_0_s1_translator:av_writedata -> new_sdram_controller_0:az_data
	wire  [21:0] new_sdram_controller_0_s1_translator_avalon_anti_slave_0_address;                               // new_sdram_controller_0_s1_translator:av_address -> new_sdram_controller_0:az_addr
	wire         new_sdram_controller_0_s1_translator_avalon_anti_slave_0_chipselect;                            // new_sdram_controller_0_s1_translator:av_chipselect -> new_sdram_controller_0:az_cs
	wire         new_sdram_controller_0_s1_translator_avalon_anti_slave_0_write;                                 // new_sdram_controller_0_s1_translator:av_write -> new_sdram_controller_0:az_wr_n
	wire         new_sdram_controller_0_s1_translator_avalon_anti_slave_0_read;                                  // new_sdram_controller_0_s1_translator:av_read -> new_sdram_controller_0:az_rd_n
	wire  [15:0] new_sdram_controller_0_s1_translator_avalon_anti_slave_0_readdata;                              // new_sdram_controller_0:za_data -> new_sdram_controller_0_s1_translator:av_readdata
	wire         new_sdram_controller_0_s1_translator_avalon_anti_slave_0_readdatavalid;                         // new_sdram_controller_0:za_valid -> new_sdram_controller_0_s1_translator:av_readdatavalid
	wire   [1:0] new_sdram_controller_0_s1_translator_avalon_anti_slave_0_byteenable;                            // new_sdram_controller_0_s1_translator:av_byteenable -> new_sdram_controller_0:az_be_n
	wire         bridge_0_avalon_master_translator_avalon_universal_master_0_waitrequest;                        // bridge_0_avalon_master_translator_avalon_universal_master_0_agent:av_waitrequest -> bridge_0_avalon_master_translator:uav_waitrequest
	wire   [1:0] bridge_0_avalon_master_translator_avalon_universal_master_0_burstcount;                         // bridge_0_avalon_master_translator:uav_burstcount -> bridge_0_avalon_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [15:0] bridge_0_avalon_master_translator_avalon_universal_master_0_writedata;                          // bridge_0_avalon_master_translator:uav_writedata -> bridge_0_avalon_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [22:0] bridge_0_avalon_master_translator_avalon_universal_master_0_address;                            // bridge_0_avalon_master_translator:uav_address -> bridge_0_avalon_master_translator_avalon_universal_master_0_agent:av_address
	wire         bridge_0_avalon_master_translator_avalon_universal_master_0_lock;                               // bridge_0_avalon_master_translator:uav_lock -> bridge_0_avalon_master_translator_avalon_universal_master_0_agent:av_lock
	wire         bridge_0_avalon_master_translator_avalon_universal_master_0_write;                              // bridge_0_avalon_master_translator:uav_write -> bridge_0_avalon_master_translator_avalon_universal_master_0_agent:av_write
	wire         bridge_0_avalon_master_translator_avalon_universal_master_0_read;                               // bridge_0_avalon_master_translator:uav_read -> bridge_0_avalon_master_translator_avalon_universal_master_0_agent:av_read
	wire  [15:0] bridge_0_avalon_master_translator_avalon_universal_master_0_readdata;                           // bridge_0_avalon_master_translator_avalon_universal_master_0_agent:av_readdata -> bridge_0_avalon_master_translator:uav_readdata
	wire         bridge_0_avalon_master_translator_avalon_universal_master_0_debugaccess;                        // bridge_0_avalon_master_translator:uav_debugaccess -> bridge_0_avalon_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [1:0] bridge_0_avalon_master_translator_avalon_universal_master_0_byteenable;                         // bridge_0_avalon_master_translator:uav_byteenable -> bridge_0_avalon_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         bridge_0_avalon_master_translator_avalon_universal_master_0_readdatavalid;                      // bridge_0_avalon_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> bridge_0_avalon_master_translator:uav_readdatavalid
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // new_sdram_controller_0_s1_translator:uav_waitrequest -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [1:0] new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;              // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> new_sdram_controller_0_s1_translator:uav_burstcount
	wire  [15:0] new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;               // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> new_sdram_controller_0_s1_translator:uav_writedata
	wire  [22:0] new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                 // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> new_sdram_controller_0_s1_translator:uav_address
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                   // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> new_sdram_controller_0_s1_translator:uav_write
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                    // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> new_sdram_controller_0_s1_translator:uav_lock
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                    // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> new_sdram_controller_0_s1_translator:uav_read
	wire  [15:0] new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                // new_sdram_controller_0_s1_translator:uav_readdata -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // new_sdram_controller_0_s1_translator:uav_readdatavalid -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> new_sdram_controller_0_s1_translator:uav_debugaccess
	wire   [1:0] new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;              // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> new_sdram_controller_0_s1_translator:uav_byteenable
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;            // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [71:0] new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;             // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;            // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [71:0] new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire  [17:0] new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;       // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [17:0] new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;        // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;       // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire         bridge_0_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket;               // bridge_0_avalon_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire         bridge_0_avalon_master_translator_avalon_universal_master_0_agent_cp_valid;                     // bridge_0_avalon_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire         bridge_0_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket;             // bridge_0_avalon_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [70:0] bridge_0_avalon_master_translator_avalon_universal_master_0_agent_cp_data;                      // bridge_0_avalon_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire         bridge_0_avalon_master_translator_avalon_universal_master_0_agent_cp_ready;                     // addr_router:sink_ready -> bridge_0_avalon_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                   // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [70:0] new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                    // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router:sink_ready -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         rst_controller_reset_out_reset;                                                                 // rst_controller:reset_out -> [addr_router:reset, bridge_0:reset, bridge_0_avalon_master_translator:reset, bridge_0_avalon_master_translator_avalon_universal_master_0_agent:reset, cmd_xbar_demux:reset, crosser:in_reset, crosser_001:out_reset, up_clocks_0:reset]
	wire         rst_controller_001_reset_out_reset;                                                             // rst_controller_001:reset_out -> [crosser:out_reset, crosser_001:in_reset, id_router:reset, new_sdram_controller_0:reset_n, new_sdram_controller_0_s1_translator:reset, new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:reset, new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset]
	wire         addr_router_src_endofpacket;                                                                    // addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire         addr_router_src_valid;                                                                          // addr_router:src_valid -> cmd_xbar_demux:sink_valid
	wire         addr_router_src_startofpacket;                                                                  // addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [70:0] addr_router_src_data;                                                                           // addr_router:src_data -> cmd_xbar_demux:sink_data
	wire   [0:0] addr_router_src_channel;                                                                        // addr_router:src_channel -> cmd_xbar_demux:sink_channel
	wire         addr_router_src_ready;                                                                          // cmd_xbar_demux:sink_ready -> addr_router:src_ready
	wire         crosser_001_out_ready;                                                                          // bridge_0_avalon_master_translator_avalon_universal_master_0_agent:rp_ready -> crosser_001:out_ready
	wire         crosser_out_ready;                                                                              // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> crosser:out_ready
	wire         id_router_src_endofpacket;                                                                      // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire         id_router_src_valid;                                                                            // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire         id_router_src_startofpacket;                                                                    // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [70:0] id_router_src_data;                                                                             // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [0:0] id_router_src_channel;                                                                          // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire         id_router_src_ready;                                                                            // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire         crosser_out_endofpacket;                                                                        // crosser:out_endofpacket -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         crosser_out_valid;                                                                              // crosser:out_valid -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         crosser_out_startofpacket;                                                                      // crosser:out_startofpacket -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [70:0] crosser_out_data;                                                                               // crosser:out_data -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire         crosser_out_channel;                                                                            // crosser:out_channel -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_src0_endofpacket;                                                                // cmd_xbar_demux:src0_endofpacket -> crosser:in_endofpacket
	wire         cmd_xbar_demux_src0_valid;                                                                      // cmd_xbar_demux:src0_valid -> crosser:in_valid
	wire         cmd_xbar_demux_src0_startofpacket;                                                              // cmd_xbar_demux:src0_startofpacket -> crosser:in_startofpacket
	wire  [70:0] cmd_xbar_demux_src0_data;                                                                       // cmd_xbar_demux:src0_data -> crosser:in_data
	wire   [0:0] cmd_xbar_demux_src0_channel;                                                                    // cmd_xbar_demux:src0_channel -> crosser:in_channel
	wire         cmd_xbar_demux_src0_ready;                                                                      // crosser:in_ready -> cmd_xbar_demux:src0_ready
	wire         crosser_001_out_endofpacket;                                                                    // crosser_001:out_endofpacket -> bridge_0_avalon_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         crosser_001_out_valid;                                                                          // crosser_001:out_valid -> bridge_0_avalon_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         crosser_001_out_startofpacket;                                                                  // crosser_001:out_startofpacket -> bridge_0_avalon_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [70:0] crosser_001_out_data;                                                                           // crosser_001:out_data -> bridge_0_avalon_master_translator_avalon_universal_master_0_agent:rp_data
	wire         crosser_001_out_channel;                                                                        // crosser_001:out_channel -> bridge_0_avalon_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_demux_src0_endofpacket;                                                                // rsp_xbar_demux:src0_endofpacket -> crosser_001:in_endofpacket
	wire         rsp_xbar_demux_src0_valid;                                                                      // rsp_xbar_demux:src0_valid -> crosser_001:in_valid
	wire         rsp_xbar_demux_src0_startofpacket;                                                              // rsp_xbar_demux:src0_startofpacket -> crosser_001:in_startofpacket
	wire  [70:0] rsp_xbar_demux_src0_data;                                                                       // rsp_xbar_demux:src0_data -> crosser_001:in_data
	wire   [0:0] rsp_xbar_demux_src0_channel;                                                                    // rsp_xbar_demux:src0_channel -> crosser_001:in_channel
	wire         rsp_xbar_demux_src0_ready;                                                                      // crosser_001:in_ready -> rsp_xbar_demux:src0_ready

	sdram_system_up_clocks_0 up_clocks_0 (
		.CLOCK_50    (clk_clk),                        //       clk_in_primary.clk
		.reset       (rst_controller_reset_out_reset), // clk_in_primary_reset.reset
		.sys_clk     (),                               //              sys_clk.clk
		.sys_reset_n (),                               //        sys_clk_reset.reset_n
		.SDRAM_CLK   (up_clocks_0_sdram_clk_clk),      //            sdram_clk.clk
		.VGA_CLK     (vga_clk_clk)                     //              vga_clk.clk
	);

	sdram_system_new_sdram_controller_0 new_sdram_controller_0 (
		.clk            (up_clocks_0_sdram_clk_clk),                                              //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),                                    // reset.reset_n
		.az_addr        (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_address),       //    s1.address
		.az_be_n        (~new_sdram_controller_0_s1_translator_avalon_anti_slave_0_byteenable),   //      .byteenable_n
		.az_cs          (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_chipselect),    //      .chipselect
		.az_data        (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.az_rd_n        (~new_sdram_controller_0_s1_translator_avalon_anti_slave_0_read),         //      .read_n
		.az_wr_n        (~new_sdram_controller_0_s1_translator_avalon_anti_slave_0_write),        //      .write_n
		.za_data        (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.za_valid       (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.za_waitrequest (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_controller_addr),                                                  //  wire.export
		.zs_ba          (sdram_controller_ba),                                                    //      .export
		.zs_cas_n       (sdram_controller_cas_n),                                                 //      .export
		.zs_cke         (sdram_controller_cke),                                                   //      .export
		.zs_cs_n        (sdram_controller_cs_n),                                                  //      .export
		.zs_dq          (sdram_controller_dq),                                                    //      .export
		.zs_dqm         (sdram_controller_dqm),                                                   //      .export
		.zs_ras_n       (sdram_controller_ras_n),                                                 //      .export
		.zs_we_n        (sdram_controller_we_n)                                                   //      .export
	);

	sdram_system_bridge_0 bridge_0 (
		.clk                (clk_clk),                            //        clock_reset.clk
		.reset              (rst_controller_reset_out_reset),     //  clock_reset_reset.reset
		.avalon_readdata    (bridge_0_avalon_master_readdata),    //      avalon_master.readdata
		.avalon_waitrequest (bridge_0_avalon_master_waitrequest), //                   .waitrequest
		.avalon_byteenable  (bridge_0_avalon_master_byteenable),  //                   .byteenable
		.avalon_read        (bridge_0_avalon_master_read),        //                   .read
		.avalon_write       (bridge_0_avalon_master_write),       //                   .write
		.avalon_writedata   (bridge_0_avalon_master_writedata),   //                   .writedata
		.avalon_address     (bridge_0_avalon_master_address),     //                   .address
		.address            (avalon_bridge_address),              // external_interface.export
		.byte_enable        (avalon_bridge_byte_enable),          //                   .export
		.read               (avalon_bridge_read),                 //                   .export
		.write              (avalon_bridge_write),                //                   .export
		.write_data         (avalon_bridge_write_data),           //                   .export
		.acknowledge        (avalon_bridge_acknowledge),          //                   .export
		.read_data          (avalon_bridge_read_data)             //                   .export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (23),
		.AV_DATA_W                   (16),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (2),
		.UAV_ADDRESS_W               (23),
		.UAV_BURSTCOUNT_W            (2),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (2),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) bridge_0_avalon_master_translator (
		.clk                      (clk_clk),                                                                   //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                            //                     reset.reset
		.uav_address              (bridge_0_avalon_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (bridge_0_avalon_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (bridge_0_avalon_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (bridge_0_avalon_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (bridge_0_avalon_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (bridge_0_avalon_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (bridge_0_avalon_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (bridge_0_avalon_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (bridge_0_avalon_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (bridge_0_avalon_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (bridge_0_avalon_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (bridge_0_avalon_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (bridge_0_avalon_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (bridge_0_avalon_master_byteenable),                                         //                          .byteenable
		.av_read                  (bridge_0_avalon_master_read),                                               //                          .read
		.av_readdata              (bridge_0_avalon_master_readdata),                                           //                          .readdata
		.av_write                 (bridge_0_avalon_master_write),                                              //                          .write
		.av_writedata             (bridge_0_avalon_master_writedata),                                          //                          .writedata
		.av_burstcount            (1'b1),                                                                      //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                      //               (terminated)
		.av_begintransfer         (1'b0),                                                                      //               (terminated)
		.av_chipselect            (1'b0),                                                                      //               (terminated)
		.av_readdatavalid         (),                                                                          //               (terminated)
		.av_lock                  (1'b0),                                                                      //               (terminated)
		.av_debugaccess           (1'b0),                                                                      //               (terminated)
		.uav_clken                (),                                                                          //               (terminated)
		.av_clken                 (1'b1),                                                                      //               (terminated)
		.uav_response             (2'b00),                                                                     //               (terminated)
		.av_response              (),                                                                          //               (terminated)
		.uav_writeresponserequest (),                                                                          //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                      //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                      //               (terminated)
		.av_writeresponsevalid    ()                                                                           //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (22),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (23),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) new_sdram_controller_0_s1_translator (
		.clk                      (up_clocks_0_sdram_clk_clk),                                                            //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                                   //                    reset.reset
		.uav_address              (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                     //              (terminated)
		.av_beginbursttransfer    (),                                                                                     //              (terminated)
		.av_burstcount            (),                                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                                     //              (terminated)
		.av_lock                  (),                                                                                     //              (terminated)
		.av_clken                 (),                                                                                     //              (terminated)
		.uav_clken                (1'b0),                                                                                 //              (terminated)
		.av_debugaccess           (),                                                                                     //              (terminated)
		.av_outputenable          (),                                                                                     //              (terminated)
		.uav_response             (),                                                                                     //              (terminated)
		.av_response              (2'b00),                                                                                //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                 //              (terminated)
		.uav_writeresponsevalid   (),                                                                                     //              (terminated)
		.av_writeresponserequest  (),                                                                                     //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                  //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (64),
		.PKT_PROTECTION_L          (62),
		.PKT_BEGIN_BURST           (57),
		.PKT_BURSTWRAP_H           (49),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BURST_SIZE_H          (52),
		.PKT_BURST_SIZE_L          (50),
		.PKT_BURST_TYPE_H          (54),
		.PKT_BURST_TYPE_L          (53),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (47),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_TRANS_EXCLUSIVE       (46),
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_SRC_ID_H              (59),
		.PKT_SRC_ID_L              (59),
		.PKT_DEST_ID_H             (60),
		.PKT_DEST_ID_L             (60),
		.PKT_THREAD_ID_H           (61),
		.PKT_THREAD_ID_L           (61),
		.PKT_CACHE_H               (68),
		.PKT_CACHE_L               (65),
		.PKT_DATA_SIDEBAND_H       (56),
		.PKT_DATA_SIDEBAND_L       (56),
		.PKT_QOS_H                 (58),
		.PKT_QOS_L                 (58),
		.PKT_ADDR_SIDEBAND_H       (55),
		.PKT_ADDR_SIDEBAND_L       (55),
		.PKT_RESPONSE_STATUS_H     (70),
		.PKT_RESPONSE_STATUS_L     (69),
		.ST_DATA_W                 (71),
		.ST_CHANNEL_W              (1),
		.AV_BURSTCOUNT_W           (2),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (1),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) bridge_0_avalon_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_clk),                                                                            //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.av_address              (bridge_0_avalon_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (bridge_0_avalon_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (bridge_0_avalon_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (bridge_0_avalon_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (bridge_0_avalon_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (bridge_0_avalon_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (bridge_0_avalon_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (bridge_0_avalon_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (bridge_0_avalon_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (bridge_0_avalon_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (bridge_0_avalon_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (bridge_0_avalon_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (bridge_0_avalon_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (bridge_0_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (bridge_0_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (bridge_0_avalon_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (crosser_001_out_valid),                                                              //        rp.valid
		.rp_data                 (crosser_001_out_data),                                                               //          .data
		.rp_channel              (crosser_001_out_channel),                                                            //          .channel
		.rp_startofpacket        (crosser_001_out_startofpacket),                                                      //          .startofpacket
		.rp_endofpacket          (crosser_001_out_endofpacket),                                                        //          .endofpacket
		.rp_ready                (crosser_001_out_ready),                                                              //          .ready
		.av_response             (),                                                                                   // (terminated)
		.av_writeresponserequest (1'b0),                                                                               // (terminated)
		.av_writeresponsevalid   ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (57),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (59),
		.PKT_SRC_ID_L              (59),
		.PKT_DEST_ID_H             (60),
		.PKT_DEST_ID_L             (60),
		.PKT_BURSTWRAP_H           (49),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (47),
		.PKT_PROTECTION_H          (64),
		.PKT_PROTECTION_L          (62),
		.PKT_RESPONSE_STATUS_H     (70),
		.PKT_RESPONSE_STATUS_L     (69),
		.PKT_BURST_SIZE_H          (52),
		.PKT_BURST_SIZE_L          (50),
		.ST_CHANNEL_W              (1),
		.ST_DATA_W                 (71),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (up_clocks_0_sdram_clk_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                             //       clk_reset.reset
		.m0_address              (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_out_ready),                                                                              //              cp.ready
		.cp_valid                (crosser_out_valid),                                                                              //                .valid
		.cp_data                 (crosser_out_data),                                                                               //                .data
		.cp_startofpacket        (crosser_out_startofpacket),                                                                      //                .startofpacket
		.cp_endofpacket          (crosser_out_endofpacket),                                                                        //                .endofpacket
		.cp_channel              (crosser_out_channel),                                                                            //                .channel
		.rf_sink_ready           (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                          //     (terminated)
		.m0_writeresponserequest (),                                                                                               //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                            //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (72),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (up_clocks_0_sdram_clk_clk),                                                                      //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                             // clk_reset.reset
		.in_data           (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                          // (terminated)
		.csr_read          (1'b0),                                                                                           // (terminated)
		.csr_write         (1'b0),                                                                                           // (terminated)
		.csr_readdata      (),                                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                           // (terminated)
		.almost_full_data  (),                                                                                               // (terminated)
		.almost_empty_data (),                                                                                               // (terminated)
		.in_empty          (1'b0),                                                                                           // (terminated)
		.out_empty         (),                                                                                               // (terminated)
		.in_error          (1'b0),                                                                                           // (terminated)
		.out_error         (),                                                                                               // (terminated)
		.in_channel        (1'b0),                                                                                           // (terminated)
		.out_channel       ()                                                                                                // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (18),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (up_clocks_0_sdram_clk_clk),                                                                //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_startofpacket  (1'b0),                                                                                     // (terminated)
		.in_endofpacket    (1'b0),                                                                                     // (terminated)
		.out_startofpacket (),                                                                                         // (terminated)
		.out_endofpacket   (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	sdram_system_addr_router addr_router (
		.sink_ready         (bridge_0_avalon_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (bridge_0_avalon_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (bridge_0_avalon_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (bridge_0_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (bridge_0_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                              //       src.ready
		.src_valid          (addr_router_src_valid),                                                              //          .valid
		.src_data           (addr_router_src_data),                                                               //          .data
		.src_channel        (addr_router_src_channel),                                                            //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                         //          .endofpacket
	);

	sdram_system_id_router id_router (
		.sink_ready         (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (up_clocks_0_sdram_clk_clk),                                                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_src_valid),                                                                  //          .valid
		.src_data           (id_router_src_data),                                                                   //          .data
		.src_channel        (id_router_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                             //          .endofpacket
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                 // reset_in0.reset
		.clk        (clk_clk),                        //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req  (),                               // (terminated)
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_001 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.clk        (up_clocks_0_sdram_clk_clk),          //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	sdram_system_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clk_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_src_ready),             //      sink.ready
		.sink_channel       (addr_router_src_channel),           //          .channel
		.sink_data          (addr_router_src_data),              //          .data
		.sink_startofpacket (addr_router_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket)    //          .endofpacket
	);

	sdram_system_cmd_xbar_demux rsp_xbar_demux (
		.clk                (up_clocks_0_sdram_clk_clk),          //       clk.clk
		.reset              (rst_controller_001_reset_out_reset), // clk_reset.reset
		.sink_ready         (id_router_src_ready),                //      sink.ready
		.sink_channel       (id_router_src_channel),              //          .channel
		.sink_data          (id_router_src_data),                 //          .data
		.sink_startofpacket (id_router_src_startofpacket),        //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),          //          .endofpacket
		.sink_valid         (id_router_src_valid),                //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),          //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),          //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),           //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),        //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket)     //          .endofpacket
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (71),
		.BITS_PER_SYMBOL     (71),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (1),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser (
		.in_clk            (clk_clk),                            //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),     //  in_clk_reset.reset
		.out_clk           (up_clocks_0_sdram_clk_clk),          //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset), // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_src0_ready),          //            in.ready
		.in_valid          (cmd_xbar_demux_src0_valid),          //              .valid
		.in_startofpacket  (cmd_xbar_demux_src0_startofpacket),  //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src0_endofpacket),    //              .endofpacket
		.in_channel        (cmd_xbar_demux_src0_channel),        //              .channel
		.in_data           (cmd_xbar_demux_src0_data),           //              .data
		.out_ready         (crosser_out_ready),                  //           out.ready
		.out_valid         (crosser_out_valid),                  //              .valid
		.out_startofpacket (crosser_out_startofpacket),          //              .startofpacket
		.out_endofpacket   (crosser_out_endofpacket),            //              .endofpacket
		.out_channel       (crosser_out_channel),                //              .channel
		.out_data          (crosser_out_data),                   //              .data
		.in_empty          (1'b0),                               //   (terminated)
		.in_error          (1'b0),                               //   (terminated)
		.out_empty         (),                                   //   (terminated)
		.out_error         ()                                    //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (71),
		.BITS_PER_SYMBOL     (71),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (1),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_001 (
		.in_clk            (up_clocks_0_sdram_clk_clk),          //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset), //  in_clk_reset.reset
		.out_clk           (clk_clk),                            //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),     // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_src0_ready),          //            in.ready
		.in_valid          (rsp_xbar_demux_src0_valid),          //              .valid
		.in_startofpacket  (rsp_xbar_demux_src0_startofpacket),  //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_src0_endofpacket),    //              .endofpacket
		.in_channel        (rsp_xbar_demux_src0_channel),        //              .channel
		.in_data           (rsp_xbar_demux_src0_data),           //              .data
		.out_ready         (crosser_001_out_ready),              //           out.ready
		.out_valid         (crosser_001_out_valid),              //              .valid
		.out_startofpacket (crosser_001_out_startofpacket),      //              .startofpacket
		.out_endofpacket   (crosser_001_out_endofpacket),        //              .endofpacket
		.out_channel       (crosser_001_out_channel),            //              .channel
		.out_data          (crosser_001_out_data),               //              .data
		.in_empty          (1'b0),                               //   (terminated)
		.in_error          (1'b0),                               //   (terminated)
		.out_empty         (),                                   //   (terminated)
		.out_error         ()                                    //   (terminated)
	);

endmodule
