module gpu(
    input CLOCK_50,
    input reset,
    input VGA_CLK,
    output wire [3:0] VGA_R,
    output wire [3:0] VGA_G,
    output wire [3:0] VGA_B,
    output wire VGA_HS,
    output wire VGA_VS
);

// Size of the text display.
parameter text_display_rows = 5'd24;
parameter text_display_columns = 7'd80;
parameter display_width_pixels = 10'd640;
parameter display_height_pixels = 9'd480;

parameter character_cell_width = display_width_pixels / text_display_columns;
parameter character_cell_height = display_height_pixels / text_display_rows;

integer i;
integer j;

// Buffer holding the text that is being displayed on-screen. Each cell in the 2-D array is a byte (8 bits) storing an ASCII character.
reg[7:0] text_buffer[text_display_rows - 1:0][text_display_columns - 1:0];

// Create a VGA controller with 25 MHz pixel clock.
wire blanking;
wire[9:0] pixel_x;
wire[8:0] pixel_y;
vga640x480 vga(.i_clk(CLOCK_50),
               .i_pix_stb(VGA_CLK),
               .i_rst(~reset),
               .o_hs(VGA_HS),
               .o_vs(VGA_VS),
               .o_blanking(blanking),
               .o_x(pixel_x),
               .o_y(pixel_y));

// Registers for tracking the coordinates of the current pixel being drawn within the current character cell.
reg[$clog2(character_cell_width) - 1:0] character_cell_x; // Units: pixels, Range: 0 to character_cell_width - 1
reg[$clog2(character_cell_height) - 1:0] character_cell_y; // Units: pixels, Range: 0 to character_cell_height - 1
// Registers for tracking the current character cell's location.
reg[$clog2(text_display_rows) - 1:0] current_row; // Units: rows of text, Range: 0 to text_display_rows - 1
reg[$clog2(text_display_columns) - 1:0] current_column; // Units: columns of text, Range: 0 to text_display_columns - 1

// Combinational logic for rendering pixels.
wire[7:0] current_character; // The character currently being drawn.
wire current_pixel_value; // The value (on or off) of the pixel currently being rendered. Generated by the font_rom module.
assign current_character = text_buffer[current_row][current_column]; // The current character is selected from the text buffer using the row and column counters.
// If we're in VGA blanking, then switch off the VGA color pins. Otherwise, use current_pixel_value to set the VGA color pins' values.
assign VGA_R = blanking ? 4'b0000 : (current_pixel_value ? 4'b1111 : 4'b0000);
assign VGA_G = blanking ? 4'b0000 : (current_pixel_value ? 4'b1111 : 4'b0000);
assign VGA_B = blanking ? 4'b0000 : (current_pixel_value ? 4'b1111 : 4'b0000);

// Font glyph lookup table, used to render text characters by determining whether the current pixel should be black or white.
font_rom font_glyphs(.character(current_character),
                     .character_cell_x(character_cell_x),
                     .character_cell_y(character_cell_y),
                     .pixel_value(current_pixel_value));

// Sequential logic for counting pixels, rows, and columns.
always @(posedge VGA_CLK)
begin
    if (reset)
    begin
        for (i = 3; i < text_display_rows; i = i + 1)
        begin
            for (j = 0; j < text_display_columns; j = j + 1)
            begin
                text_buffer[i][j] <= 'd0;
            end
        end
        for (j = 1; j < text_display_columns - 1; j = j + 1)
            text_buffer[0][j] <= 'd65;
        text_buffer[0][0] <= 'd35;
        text_buffer[0][text_display_columns - 1] <= 'd36;
        for (j = 0; j < text_display_columns; j = j + 1)
            text_buffer[1][j] <= 'd66;
        for (j = 0; j < text_display_columns; j = j + 1)
            text_buffer[2][j] <= 'd67;
        character_cell_x <= 'h0;
        character_cell_y <= 'h0;
        current_row <= 'h0;
        current_column <= 'h0;
        $display("In reset.");
    end
    else if (~blanking)
    begin
        $display("Rendering.");
        if (current_column == text_display_columns)
        begin
            character_cell_x <= 'd0;
            current_column <= 'd0;
        end
        else
        begin
            if (character_cell_x + 'd1 == character_cell_width)
            begin
                character_cell_x <= 'd0;
                current_column <= current_column + 'd1;
            end
            else
                character_cell_x <= character_cell_x + 'd1;
        end

        if (pixel_x == 0 && pixel_y == 0)
        begin
            character_cell_y <= 'd0;
            current_row <= 'd0;
        end
        else
        begin
            if (character_cell_y == character_cell_height)
            begin
                character_cell_y <= 'd0;
                current_row <= current_row + 'd1;
            end
            else if (pixel_x == display_width_pixels)
                character_cell_y <= character_cell_y + 'd1;
        end
    end
end

endmodule
