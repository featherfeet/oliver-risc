module rom(input[31:0] address, output reg [7:0] output_byte, output done);
	assign done = (address == 32'd1866) ? 1'b1 : 1'b0;
	always @(address)
	begin
		case (address)
			32'd0:
				output_byte = 8'd0;
			32'd1:
				output_byte = 8'd0;
			32'd2:
				output_byte = 8'd0;
			32'd3:
				output_byte = 8'd0;
			32'd4:
				output_byte = 8'd0;
			32'd5:
				output_byte = 8'd0;
			32'd6:
				output_byte = 8'd0;
			32'd7:
				output_byte = 8'd0;
			32'd8:
				output_byte = 8'd0;
			32'd9:
				output_byte = 8'd0;
			32'd10:
				output_byte = 8'd0;
			32'd11:
				output_byte = 8'd0;
			32'd12:
				output_byte = 8'd0;
			32'd13:
				output_byte = 8'd0;
			32'd14:
				output_byte = 8'd0;
			32'd15:
				output_byte = 8'd0;
			32'd16:
				output_byte = 8'd0;
			32'd17:
				output_byte = 8'd0;
			32'd18:
				output_byte = 8'd0;
			32'd19:
				output_byte = 8'd0;
			32'd20:
				output_byte = 8'd0;
			32'd21:
				output_byte = 8'd0;
			32'd22:
				output_byte = 8'd0;
			32'd23:
				output_byte = 8'd0;
			32'd24:
				output_byte = 8'd0;
			32'd25:
				output_byte = 8'd0;
			32'd26:
				output_byte = 8'd0;
			32'd27:
				output_byte = 8'd0;
			32'd28:
				output_byte = 8'd0;
			32'd29:
				output_byte = 8'd0;
			32'd30:
				output_byte = 8'd0;
			32'd31:
				output_byte = 8'd0;
			32'd32:
				output_byte = 8'd0;
			32'd33:
				output_byte = 8'd0;
			32'd34:
				output_byte = 8'd0;
			32'd35:
				output_byte = 8'd0;
			32'd36:
				output_byte = 8'd0;
			32'd37:
				output_byte = 8'd0;
			32'd38:
				output_byte = 8'd0;
			32'd39:
				output_byte = 8'd0;
			32'd40:
				output_byte = 8'd0;
			32'd41:
				output_byte = 8'd0;
			32'd42:
				output_byte = 8'd0;
			32'd43:
				output_byte = 8'd0;
			32'd44:
				output_byte = 8'd0;
			32'd45:
				output_byte = 8'd0;
			32'd46:
				output_byte = 8'd0;
			32'd47:
				output_byte = 8'd0;
			32'd48:
				output_byte = 8'd14;
			32'd49:
				output_byte = 8'd20;
			32'd50:
				output_byte = 8'd4;
			32'd51:
				output_byte = 8'd0;
			32'd52:
				output_byte = 8'd0;
			32'd53:
				output_byte = 8'd0;
			32'd54:
				output_byte = 8'd1;
			32'd55:
				output_byte = 8'd0;
			32'd56:
				output_byte = 8'd0;
			32'd57:
				output_byte = 8'd0;
			32'd58:
				output_byte = 8'd2;
			32'd59:
				output_byte = 8'd1;
			32'd60:
				output_byte = 8'd0;
			32'd61:
				output_byte = 8'd0;
			32'd62:
				output_byte = 8'd0;
			32'd63:
				output_byte = 8'd8;
			32'd64:
				output_byte = 8'd0;
			32'd65:
				output_byte = 8'd0;
			32'd66:
				output_byte = 8'd0;
			32'd67:
				output_byte = 8'd20;
			32'd68:
				output_byte = 8'd0;
			32'd69:
				output_byte = 8'd0;
			32'd70:
				output_byte = 8'd0;
			32'd71:
				output_byte = 8'd0;
			32'd72:
				output_byte = 8'd1;
			32'd73:
				output_byte = 8'd0;
			32'd74:
				output_byte = 8'd0;
			32'd75:
				output_byte = 8'd0;
			32'd76:
				output_byte = 8'd2;
			32'd77:
				output_byte = 8'd1;
			32'd78:
				output_byte = 8'd0;
			32'd79:
				output_byte = 8'd0;
			32'd80:
				output_byte = 8'd0;
			32'd81:
				output_byte = 8'd12;
			32'd82:
				output_byte = 8'd0;
			32'd83:
				output_byte = 8'd0;
			32'd84:
				output_byte = 8'd0;
			32'd85:
				output_byte = 8'd20;
			32'd86:
				output_byte = 8'd2;
			32'd87:
				output_byte = 8'd0;
			32'd88:
				output_byte = 8'd0;
			32'd89:
				output_byte = 8'd0;
			32'd90:
				output_byte = 8'd1;
			32'd91:
				output_byte = 8'd0;
			32'd92:
				output_byte = 8'd0;
			32'd93:
				output_byte = 8'd0;
			32'd94:
				output_byte = 8'd2;
			32'd95:
				output_byte = 8'd1;
			32'd96:
				output_byte = 8'd0;
			32'd97:
				output_byte = 8'd0;
			32'd98:
				output_byte = 8'd0;
			32'd99:
				output_byte = 8'd16;
			32'd100:
				output_byte = 8'd0;
			32'd101:
				output_byte = 8'd0;
			32'd102:
				output_byte = 8'd0;
			32'd103:
				output_byte = 8'd20;
			32'd104:
				output_byte = 8'd80;
			32'd105:
				output_byte = 8'd0;
			32'd106:
				output_byte = 8'd0;
			32'd107:
				output_byte = 8'd0;
			32'd108:
				output_byte = 8'd1;
			32'd109:
				output_byte = 8'd0;
			32'd110:
				output_byte = 8'd0;
			32'd111:
				output_byte = 8'd0;
			32'd112:
				output_byte = 8'd2;
			32'd113:
				output_byte = 8'd1;
			32'd114:
				output_byte = 8'd0;
			32'd115:
				output_byte = 8'd0;
			32'd116:
				output_byte = 8'd0;
			32'd117:
				output_byte = 8'd20;
			32'd118:
				output_byte = 8'd0;
			32'd119:
				output_byte = 8'd0;
			32'd120:
				output_byte = 8'd0;
			32'd121:
				output_byte = 8'd20;
			32'd122:
				output_byte = 8'd2;
			32'd123:
				output_byte = 8'd0;
			32'd124:
				output_byte = 8'd0;
			32'd125:
				output_byte = 8'd0;
			32'd126:
				output_byte = 8'd1;
			32'd127:
				output_byte = 8'd0;
			32'd128:
				output_byte = 8'd0;
			32'd129:
				output_byte = 8'd0;
			32'd130:
				output_byte = 8'd2;
			32'd131:
				output_byte = 8'd1;
			32'd132:
				output_byte = 8'd0;
			32'd133:
				output_byte = 8'd0;
			32'd134:
				output_byte = 8'd0;
			32'd135:
				output_byte = 8'd24;
			32'd136:
				output_byte = 8'd0;
			32'd137:
				output_byte = 8'd0;
			32'd138:
				output_byte = 8'd0;
			32'd139:
				output_byte = 8'd20;
			32'd140:
				output_byte = 8'd0;
			32'd141:
				output_byte = 8'd0;
			32'd142:
				output_byte = 8'd0;
			32'd143:
				output_byte = 8'd0;
			32'd144:
				output_byte = 8'd1;
			32'd145:
				output_byte = 8'd0;
			32'd146:
				output_byte = 8'd0;
			32'd147:
				output_byte = 8'd0;
			32'd148:
				output_byte = 8'd2;
			32'd149:
				output_byte = 8'd1;
			32'd150:
				output_byte = 8'd0;
			32'd151:
				output_byte = 8'd0;
			32'd152:
				output_byte = 8'd0;
			32'd153:
				output_byte = 8'd28;
			32'd154:
				output_byte = 8'd0;
			32'd155:
				output_byte = 8'd0;
			32'd156:
				output_byte = 8'd0;
			32'd157:
				output_byte = 8'd20;
			32'd158:
				output_byte = 8'd0;
			32'd159:
				output_byte = 8'd0;
			32'd160:
				output_byte = 8'd0;
			32'd161:
				output_byte = 8'd0;
			32'd162:
				output_byte = 8'd1;
			32'd163:
				output_byte = 8'd0;
			32'd164:
				output_byte = 8'd0;
			32'd165:
				output_byte = 8'd0;
			32'd166:
				output_byte = 8'd2;
			32'd167:
				output_byte = 8'd1;
			32'd168:
				output_byte = 8'd0;
			32'd169:
				output_byte = 8'd0;
			32'd170:
				output_byte = 8'd0;
			32'd171:
				output_byte = 8'd32;
			32'd172:
				output_byte = 8'd0;
			32'd173:
				output_byte = 8'd0;
			32'd174:
				output_byte = 8'd0;
			32'd175:
				output_byte = 8'd20;
			32'd176:
				output_byte = 8'd0;
			32'd177:
				output_byte = 8'd0;
			32'd178:
				output_byte = 8'd0;
			32'd179:
				output_byte = 8'd0;
			32'd180:
				output_byte = 8'd1;
			32'd181:
				output_byte = 8'd0;
			32'd182:
				output_byte = 8'd0;
			32'd183:
				output_byte = 8'd0;
			32'd184:
				output_byte = 8'd1;
			32'd185:
				output_byte = 8'd12;
			32'd186:
				output_byte = 8'd0;
			32'd187:
				output_byte = 8'd0;
			32'd188:
				output_byte = 8'd0;
			32'd189:
				output_byte = 8'd2;
			32'd190:
				output_byte = 8'd0;
			32'd191:
				output_byte = 8'd0;
			32'd192:
				output_byte = 8'd0;
			32'd193:
				output_byte = 8'd3;
			32'd194:
				output_byte = 8'd1;
			32'd195:
				output_byte = 8'd0;
			32'd196:
				output_byte = 8'd0;
			32'd197:
				output_byte = 8'd0;
			32'd198:
				output_byte = 8'd2;
			32'd199:
				output_byte = 8'd0;
			32'd200:
				output_byte = 8'd0;
			32'd201:
				output_byte = 8'd0;
			32'd202:
				output_byte = 8'd7;
			32'd203:
				output_byte = 8'd1;
			32'd204:
				output_byte = 8'd0;
			32'd205:
				output_byte = 8'd0;
			32'd206:
				output_byte = 8'd0;
			32'd207:
				output_byte = 8'd3;
			32'd208:
				output_byte = 8'd0;
			32'd209:
				output_byte = 8'd0;
			32'd210:
				output_byte = 8'd0;
			32'd211:
				output_byte = 8'd20;
			32'd212:
				output_byte = 8'd0;
			32'd213:
				output_byte = 8'd0;
			32'd214:
				output_byte = 8'd0;
			32'd215:
				output_byte = 8'd0;
			32'd216:
				output_byte = 8'd1;
			32'd217:
				output_byte = 8'd0;
			32'd218:
				output_byte = 8'd0;
			32'd219:
				output_byte = 8'd0;
			32'd220:
				output_byte = 8'd1;
			32'd221:
				output_byte = 8'd8;
			32'd222:
				output_byte = 8'd0;
			32'd223:
				output_byte = 8'd0;
			32'd224:
				output_byte = 8'd0;
			32'd225:
				output_byte = 8'd2;
			32'd226:
				output_byte = 8'd0;
			32'd227:
				output_byte = 8'd0;
			32'd228:
				output_byte = 8'd0;
			32'd229:
				output_byte = 8'd3;
			32'd230:
				output_byte = 8'd1;
			32'd231:
				output_byte = 8'd0;
			32'd232:
				output_byte = 8'd0;
			32'd233:
				output_byte = 8'd0;
			32'd234:
				output_byte = 8'd2;
			32'd235:
				output_byte = 8'd0;
			32'd236:
				output_byte = 8'd0;
			32'd237:
				output_byte = 8'd0;
			32'd238:
				output_byte = 8'd8;
			32'd239:
				output_byte = 8'd3;
			32'd240:
				output_byte = 8'd0;
			32'd241:
				output_byte = 8'd0;
			32'd242:
				output_byte = 8'd0;
			32'd243:
				output_byte = 8'd1;
			32'd244:
				output_byte = 8'd0;
			32'd245:
				output_byte = 8'd0;
			32'd246:
				output_byte = 8'd0;
			32'd247:
				output_byte = 8'd10;
			32'd248:
				output_byte = 8'd17;
			32'd249:
				output_byte = 8'd7;
			32'd250:
				output_byte = 8'd0;
			32'd251:
				output_byte = 8'd0;
			32'd252:
				output_byte = 8'd0;
			32'd253:
				output_byte = 8'd0;
			32'd254:
				output_byte = 8'd0;
			32'd255:
				output_byte = 8'd0;
			32'd256:
				output_byte = 8'd11;
			32'd257:
				output_byte = 8'd17;
			32'd258:
				output_byte = 8'd7;
			32'd259:
				output_byte = 8'd0;
			32'd260:
				output_byte = 8'd0;
			32'd261:
				output_byte = 8'd0;
			32'd262:
				output_byte = 8'd0;
			32'd263:
				output_byte = 8'd0;
			32'd264:
				output_byte = 8'd0;
			32'd265:
				output_byte = 8'd20;
			32'd266:
				output_byte = 8'd0;
			32'd267:
				output_byte = 8'd0;
			32'd268:
				output_byte = 8'd0;
			32'd269:
				output_byte = 8'd0;
			32'd270:
				output_byte = 8'd1;
			32'd271:
				output_byte = 8'd0;
			32'd272:
				output_byte = 8'd0;
			32'd273:
				output_byte = 8'd0;
			32'd274:
				output_byte = 8'd20;
			32'd275:
				output_byte = 8'd2;
			32'd276:
				output_byte = 8'd0;
			32'd277:
				output_byte = 8'd0;
			32'd278:
				output_byte = 8'd0;
			32'd279:
				output_byte = 8'd2;
			32'd280:
				output_byte = 8'd0;
			32'd281:
				output_byte = 8'd0;
			32'd282:
				output_byte = 8'd0;
			32'd283:
				output_byte = 8'd3;
			32'd284:
				output_byte = 8'd1;
			32'd285:
				output_byte = 8'd0;
			32'd286:
				output_byte = 8'd0;
			32'd287:
				output_byte = 8'd0;
			32'd288:
				output_byte = 8'd2;
			32'd289:
				output_byte = 8'd0;
			32'd290:
				output_byte = 8'd0;
			32'd291:
				output_byte = 8'd0;
			32'd292:
				output_byte = 8'd2;
			32'd293:
				output_byte = 8'd1;
			32'd294:
				output_byte = 8'd0;
			32'd295:
				output_byte = 8'd0;
			32'd296:
				output_byte = 8'd0;
			32'd297:
				output_byte = 8'd24;
			32'd298:
				output_byte = 8'd0;
			32'd299:
				output_byte = 8'd0;
			32'd300:
				output_byte = 8'd0;
			32'd301:
				output_byte = 8'd20;
			32'd302:
				output_byte = 8'd0;
			32'd303:
				output_byte = 8'd0;
			32'd304:
				output_byte = 8'd0;
			32'd305:
				output_byte = 8'd0;
			32'd306:
				output_byte = 8'd1;
			32'd307:
				output_byte = 8'd0;
			32'd308:
				output_byte = 8'd0;
			32'd309:
				output_byte = 8'd0;
			32'd310:
				output_byte = 8'd20;
			32'd311:
				output_byte = 8'd1;
			32'd312:
				output_byte = 8'd0;
			32'd313:
				output_byte = 8'd0;
			32'd314:
				output_byte = 8'd0;
			32'd315:
				output_byte = 8'd2;
			32'd316:
				output_byte = 8'd0;
			32'd317:
				output_byte = 8'd0;
			32'd318:
				output_byte = 8'd0;
			32'd319:
				output_byte = 8'd3;
			32'd320:
				output_byte = 8'd1;
			32'd321:
				output_byte = 8'd0;
			32'd322:
				output_byte = 8'd0;
			32'd323:
				output_byte = 8'd0;
			32'd324:
				output_byte = 8'd2;
			32'd325:
				output_byte = 8'd0;
			32'd326:
				output_byte = 8'd0;
			32'd327:
				output_byte = 8'd0;
			32'd328:
				output_byte = 8'd2;
			32'd329:
				output_byte = 8'd1;
			32'd330:
				output_byte = 8'd0;
			32'd331:
				output_byte = 8'd0;
			32'd332:
				output_byte = 8'd0;
			32'd333:
				output_byte = 8'd32;
			32'd334:
				output_byte = 8'd0;
			32'd335:
				output_byte = 8'd0;
			32'd336:
				output_byte = 8'd0;
			32'd337:
				output_byte = 8'd20;
			32'd338:
				output_byte = 8'd0;
			32'd339:
				output_byte = 8'd0;
			32'd340:
				output_byte = 8'd0;
			32'd341:
				output_byte = 8'd0;
			32'd342:
				output_byte = 8'd1;
			32'd343:
				output_byte = 8'd0;
			32'd344:
				output_byte = 8'd0;
			32'd345:
				output_byte = 8'd0;
			32'd346:
				output_byte = 8'd1;
			32'd347:
				output_byte = 8'd24;
			32'd348:
				output_byte = 8'd0;
			32'd349:
				output_byte = 8'd0;
			32'd350:
				output_byte = 8'd0;
			32'd351:
				output_byte = 8'd2;
			32'd352:
				output_byte = 8'd0;
			32'd353:
				output_byte = 8'd0;
			32'd354:
				output_byte = 8'd0;
			32'd355:
				output_byte = 8'd3;
			32'd356:
				output_byte = 8'd1;
			32'd357:
				output_byte = 8'd0;
			32'd358:
				output_byte = 8'd0;
			32'd359:
				output_byte = 8'd0;
			32'd360:
				output_byte = 8'd2;
			32'd361:
				output_byte = 8'd0;
			32'd362:
				output_byte = 8'd0;
			32'd363:
				output_byte = 8'd0;
			32'd364:
				output_byte = 8'd7;
			32'd365:
				output_byte = 8'd1;
			32'd366:
				output_byte = 8'd0;
			32'd367:
				output_byte = 8'd0;
			32'd368:
				output_byte = 8'd0;
			32'd369:
				output_byte = 8'd3;
			32'd370:
				output_byte = 8'd0;
			32'd371:
				output_byte = 8'd0;
			32'd372:
				output_byte = 8'd0;
			32'd373:
				output_byte = 8'd20;
			32'd374:
				output_byte = 8'd0;
			32'd375:
				output_byte = 8'd0;
			32'd376:
				output_byte = 8'd0;
			32'd377:
				output_byte = 8'd0;
			32'd378:
				output_byte = 8'd1;
			32'd379:
				output_byte = 8'd0;
			32'd380:
				output_byte = 8'd0;
			32'd381:
				output_byte = 8'd0;
			32'd382:
				output_byte = 8'd1;
			32'd383:
				output_byte = 8'd16;
			32'd384:
				output_byte = 8'd0;
			32'd385:
				output_byte = 8'd0;
			32'd386:
				output_byte = 8'd0;
			32'd387:
				output_byte = 8'd2;
			32'd388:
				output_byte = 8'd0;
			32'd389:
				output_byte = 8'd0;
			32'd390:
				output_byte = 8'd0;
			32'd391:
				output_byte = 8'd3;
			32'd392:
				output_byte = 8'd1;
			32'd393:
				output_byte = 8'd0;
			32'd394:
				output_byte = 8'd0;
			32'd395:
				output_byte = 8'd0;
			32'd396:
				output_byte = 8'd2;
			32'd397:
				output_byte = 8'd0;
			32'd398:
				output_byte = 8'd0;
			32'd399:
				output_byte = 8'd0;
			32'd400:
				output_byte = 8'd8;
			32'd401:
				output_byte = 8'd3;
			32'd402:
				output_byte = 8'd0;
			32'd403:
				output_byte = 8'd0;
			32'd404:
				output_byte = 8'd0;
			32'd405:
				output_byte = 8'd1;
			32'd406:
				output_byte = 8'd0;
			32'd407:
				output_byte = 8'd0;
			32'd408:
				output_byte = 8'd0;
			32'd409:
				output_byte = 8'd10;
			32'd410:
				output_byte = 8'd253;
			32'd411:
				output_byte = 8'd2;
			32'd412:
				output_byte = 8'd0;
			32'd413:
				output_byte = 8'd0;
			32'd414:
				output_byte = 8'd0;
			32'd415:
				output_byte = 8'd0;
			32'd416:
				output_byte = 8'd0;
			32'd417:
				output_byte = 8'd0;
			32'd418:
				output_byte = 8'd11;
			32'd419:
				output_byte = 8'd253;
			32'd420:
				output_byte = 8'd2;
			32'd421:
				output_byte = 8'd0;
			32'd422:
				output_byte = 8'd0;
			32'd423:
				output_byte = 8'd0;
			32'd424:
				output_byte = 8'd0;
			32'd425:
				output_byte = 8'd0;
			32'd426:
				output_byte = 8'd0;
			32'd427:
				output_byte = 8'd20;
			32'd428:
				output_byte = 8'd0;
			32'd429:
				output_byte = 8'd0;
			32'd430:
				output_byte = 8'd0;
			32'd431:
				output_byte = 8'd0;
			32'd432:
				output_byte = 8'd1;
			32'd433:
				output_byte = 8'd0;
			32'd434:
				output_byte = 8'd0;
			32'd435:
				output_byte = 8'd0;
			32'd436:
				output_byte = 8'd1;
			32'd437:
				output_byte = 8'd16;
			32'd438:
				output_byte = 8'd0;
			32'd439:
				output_byte = 8'd0;
			32'd440:
				output_byte = 8'd0;
			32'd441:
				output_byte = 8'd2;
			32'd442:
				output_byte = 8'd0;
			32'd443:
				output_byte = 8'd0;
			32'd444:
				output_byte = 8'd0;
			32'd445:
				output_byte = 8'd3;
			32'd446:
				output_byte = 8'd1;
			32'd447:
				output_byte = 8'd0;
			32'd448:
				output_byte = 8'd0;
			32'd449:
				output_byte = 8'd0;
			32'd450:
				output_byte = 8'd2;
			32'd451:
				output_byte = 8'd0;
			32'd452:
				output_byte = 8'd0;
			32'd453:
				output_byte = 8'd0;
			32'd454:
				output_byte = 8'd1;
			32'd455:
				output_byte = 8'd24;
			32'd456:
				output_byte = 8'd0;
			32'd457:
				output_byte = 8'd0;
			32'd458:
				output_byte = 8'd0;
			32'd459:
				output_byte = 8'd2;
			32'd460:
				output_byte = 8'd0;
			32'd461:
				output_byte = 8'd0;
			32'd462:
				output_byte = 8'd0;
			32'd463:
				output_byte = 8'd22;
			32'd464:
				output_byte = 8'd1;
			32'd465:
				output_byte = 8'd0;
			32'd466:
				output_byte = 8'd0;
			32'd467:
				output_byte = 8'd0;
			32'd468:
				output_byte = 8'd2;
			32'd469:
				output_byte = 8'd0;
			32'd470:
				output_byte = 8'd0;
			32'd471:
				output_byte = 8'd0;
			32'd472:
				output_byte = 8'd7;
			32'd473:
				output_byte = 8'd2;
			32'd474:
				output_byte = 8'd0;
			32'd475:
				output_byte = 8'd0;
			32'd476:
				output_byte = 8'd0;
			32'd477:
				output_byte = 8'd1;
			32'd478:
				output_byte = 8'd0;
			32'd479:
				output_byte = 8'd0;
			32'd480:
				output_byte = 8'd0;
			32'd481:
				output_byte = 8'd2;
			32'd482:
				output_byte = 8'd1;
			32'd483:
				output_byte = 8'd0;
			32'd484:
				output_byte = 8'd0;
			32'd485:
				output_byte = 8'd0;
			32'd486:
				output_byte = 8'd28;
			32'd487:
				output_byte = 8'd0;
			32'd488:
				output_byte = 8'd0;
			32'd489:
				output_byte = 8'd0;
			32'd490:
				output_byte = 8'd20;
			32'd491:
				output_byte = 8'd0;
			32'd492:
				output_byte = 8'd0;
			32'd493:
				output_byte = 8'd0;
			32'd494:
				output_byte = 8'd0;
			32'd495:
				output_byte = 8'd1;
			32'd496:
				output_byte = 8'd0;
			32'd497:
				output_byte = 8'd0;
			32'd498:
				output_byte = 8'd0;
			32'd499:
				output_byte = 8'd1;
			32'd500:
				output_byte = 8'd28;
			32'd501:
				output_byte = 8'd0;
			32'd502:
				output_byte = 8'd0;
			32'd503:
				output_byte = 8'd0;
			32'd504:
				output_byte = 8'd2;
			32'd505:
				output_byte = 8'd0;
			32'd506:
				output_byte = 8'd0;
			32'd507:
				output_byte = 8'd0;
			32'd508:
				output_byte = 8'd3;
			32'd509:
				output_byte = 8'd1;
			32'd510:
				output_byte = 8'd0;
			32'd511:
				output_byte = 8'd0;
			32'd512:
				output_byte = 8'd0;
			32'd513:
				output_byte = 8'd2;
			32'd514:
				output_byte = 8'd0;
			32'd515:
				output_byte = 8'd0;
			32'd516:
				output_byte = 8'd0;
			32'd517:
				output_byte = 8'd7;
			32'd518:
				output_byte = 8'd1;
			32'd519:
				output_byte = 8'd0;
			32'd520:
				output_byte = 8'd0;
			32'd521:
				output_byte = 8'd0;
			32'd522:
				output_byte = 8'd3;
			32'd523:
				output_byte = 8'd0;
			32'd524:
				output_byte = 8'd0;
			32'd525:
				output_byte = 8'd0;
			32'd526:
				output_byte = 8'd20;
			32'd527:
				output_byte = 8'd0;
			32'd528:
				output_byte = 8'd0;
			32'd529:
				output_byte = 8'd0;
			32'd530:
				output_byte = 8'd0;
			32'd531:
				output_byte = 8'd1;
			32'd532:
				output_byte = 8'd0;
			32'd533:
				output_byte = 8'd0;
			32'd534:
				output_byte = 8'd0;
			32'd535:
				output_byte = 8'd20;
			32'd536:
				output_byte = 8'd0;
			32'd537:
				output_byte = 8'd0;
			32'd538:
				output_byte = 8'd0;
			32'd539:
				output_byte = 8'd0;
			32'd540:
				output_byte = 8'd2;
			32'd541:
				output_byte = 8'd0;
			32'd542:
				output_byte = 8'd0;
			32'd543:
				output_byte = 8'd0;
			32'd544:
				output_byte = 8'd3;
			32'd545:
				output_byte = 8'd1;
			32'd546:
				output_byte = 8'd0;
			32'd547:
				output_byte = 8'd0;
			32'd548:
				output_byte = 8'd0;
			32'd549:
				output_byte = 8'd2;
			32'd550:
				output_byte = 8'd0;
			32'd551:
				output_byte = 8'd0;
			32'd552:
				output_byte = 8'd0;
			32'd553:
				output_byte = 8'd8;
			32'd554:
				output_byte = 8'd3;
			32'd555:
				output_byte = 8'd0;
			32'd556:
				output_byte = 8'd0;
			32'd557:
				output_byte = 8'd0;
			32'd558:
				output_byte = 8'd1;
			32'd559:
				output_byte = 8'd0;
			32'd560:
				output_byte = 8'd0;
			32'd561:
				output_byte = 8'd0;
			32'd562:
				output_byte = 8'd9;
			32'd563:
				output_byte = 8'd91;
			32'd564:
				output_byte = 8'd2;
			32'd565:
				output_byte = 8'd0;
			32'd566:
				output_byte = 8'd0;
			32'd567:
				output_byte = 8'd0;
			32'd568:
				output_byte = 8'd0;
			32'd569:
				output_byte = 8'd0;
			32'd570:
				output_byte = 8'd0;
			32'd571:
				output_byte = 8'd11;
			32'd572:
				output_byte = 8'd91;
			32'd573:
				output_byte = 8'd2;
			32'd574:
				output_byte = 8'd0;
			32'd575:
				output_byte = 8'd0;
			32'd576:
				output_byte = 8'd0;
			32'd577:
				output_byte = 8'd0;
			32'd578:
				output_byte = 8'd0;
			32'd579:
				output_byte = 8'd0;
			32'd580:
				output_byte = 8'd20;
			32'd581:
				output_byte = 8'd0;
			32'd582:
				output_byte = 8'd0;
			32'd583:
				output_byte = 8'd0;
			32'd584:
				output_byte = 8'd0;
			32'd585:
				output_byte = 8'd1;
			32'd586:
				output_byte = 8'd0;
			32'd587:
				output_byte = 8'd0;
			32'd588:
				output_byte = 8'd0;
			32'd589:
				output_byte = 8'd1;
			32'd590:
				output_byte = 8'd16;
			32'd591:
				output_byte = 8'd0;
			32'd592:
				output_byte = 8'd0;
			32'd593:
				output_byte = 8'd0;
			32'd594:
				output_byte = 8'd2;
			32'd595:
				output_byte = 8'd0;
			32'd596:
				output_byte = 8'd0;
			32'd597:
				output_byte = 8'd0;
			32'd598:
				output_byte = 8'd3;
			32'd599:
				output_byte = 8'd1;
			32'd600:
				output_byte = 8'd0;
			32'd601:
				output_byte = 8'd0;
			32'd602:
				output_byte = 8'd0;
			32'd603:
				output_byte = 8'd2;
			32'd604:
				output_byte = 8'd0;
			32'd605:
				output_byte = 8'd0;
			32'd606:
				output_byte = 8'd0;
			32'd607:
				output_byte = 8'd2;
			32'd608:
				output_byte = 8'd1;
			32'd609:
				output_byte = 8'd0;
			32'd610:
				output_byte = 8'd0;
			32'd611:
				output_byte = 8'd0;
			32'd612:
				output_byte = 8'd24;
			32'd613:
				output_byte = 8'd0;
			32'd614:
				output_byte = 8'd0;
			32'd615:
				output_byte = 8'd0;
			32'd616:
				output_byte = 8'd20;
			32'd617:
				output_byte = 8'd0;
			32'd618:
				output_byte = 8'd0;
			32'd619:
				output_byte = 8'd0;
			32'd620:
				output_byte = 8'd0;
			32'd621:
				output_byte = 8'd1;
			32'd622:
				output_byte = 8'd0;
			32'd623:
				output_byte = 8'd0;
			32'd624:
				output_byte = 8'd0;
			32'd625:
				output_byte = 8'd20;
			32'd626:
				output_byte = 8'd0;
			32'd627:
				output_byte = 8'd0;
			32'd628:
				output_byte = 8'd0;
			32'd629:
				output_byte = 8'd0;
			32'd630:
				output_byte = 8'd2;
			32'd631:
				output_byte = 8'd0;
			32'd632:
				output_byte = 8'd0;
			32'd633:
				output_byte = 8'd0;
			32'd634:
				output_byte = 8'd3;
			32'd635:
				output_byte = 8'd1;
			32'd636:
				output_byte = 8'd0;
			32'd637:
				output_byte = 8'd0;
			32'd638:
				output_byte = 8'd0;
			32'd639:
				output_byte = 8'd2;
			32'd640:
				output_byte = 8'd0;
			32'd641:
				output_byte = 8'd0;
			32'd642:
				output_byte = 8'd0;
			32'd643:
				output_byte = 8'd2;
			32'd644:
				output_byte = 8'd1;
			32'd645:
				output_byte = 8'd0;
			32'd646:
				output_byte = 8'd0;
			32'd647:
				output_byte = 8'd0;
			32'd648:
				output_byte = 8'd32;
			32'd649:
				output_byte = 8'd0;
			32'd650:
				output_byte = 8'd0;
			32'd651:
				output_byte = 8'd0;
			32'd652:
				output_byte = 8'd20;
			32'd653:
				output_byte = 8'd0;
			32'd654:
				output_byte = 8'd0;
			32'd655:
				output_byte = 8'd0;
			32'd656:
				output_byte = 8'd0;
			32'd657:
				output_byte = 8'd1;
			32'd658:
				output_byte = 8'd0;
			32'd659:
				output_byte = 8'd0;
			32'd660:
				output_byte = 8'd0;
			32'd661:
				output_byte = 8'd1;
			32'd662:
				output_byte = 8'd28;
			32'd663:
				output_byte = 8'd0;
			32'd664:
				output_byte = 8'd0;
			32'd665:
				output_byte = 8'd0;
			32'd666:
				output_byte = 8'd2;
			32'd667:
				output_byte = 8'd0;
			32'd668:
				output_byte = 8'd0;
			32'd669:
				output_byte = 8'd0;
			32'd670:
				output_byte = 8'd3;
			32'd671:
				output_byte = 8'd1;
			32'd672:
				output_byte = 8'd0;
			32'd673:
				output_byte = 8'd0;
			32'd674:
				output_byte = 8'd0;
			32'd675:
				output_byte = 8'd2;
			32'd676:
				output_byte = 8'd0;
			32'd677:
				output_byte = 8'd0;
			32'd678:
				output_byte = 8'd0;
			32'd679:
				output_byte = 8'd7;
			32'd680:
				output_byte = 8'd1;
			32'd681:
				output_byte = 8'd0;
			32'd682:
				output_byte = 8'd0;
			32'd683:
				output_byte = 8'd0;
			32'd684:
				output_byte = 8'd3;
			32'd685:
				output_byte = 8'd0;
			32'd686:
				output_byte = 8'd0;
			32'd687:
				output_byte = 8'd0;
			32'd688:
				output_byte = 8'd20;
			32'd689:
				output_byte = 8'd0;
			32'd690:
				output_byte = 8'd0;
			32'd691:
				output_byte = 8'd0;
			32'd692:
				output_byte = 8'd0;
			32'd693:
				output_byte = 8'd1;
			32'd694:
				output_byte = 8'd0;
			32'd695:
				output_byte = 8'd0;
			32'd696:
				output_byte = 8'd0;
			32'd697:
				output_byte = 8'd20;
			32'd698:
				output_byte = 8'd0;
			32'd699:
				output_byte = 8'd0;
			32'd700:
				output_byte = 8'd0;
			32'd701:
				output_byte = 8'd0;
			32'd702:
				output_byte = 8'd2;
			32'd703:
				output_byte = 8'd0;
			32'd704:
				output_byte = 8'd0;
			32'd705:
				output_byte = 8'd0;
			32'd706:
				output_byte = 8'd3;
			32'd707:
				output_byte = 8'd1;
			32'd708:
				output_byte = 8'd0;
			32'd709:
				output_byte = 8'd0;
			32'd710:
				output_byte = 8'd0;
			32'd711:
				output_byte = 8'd2;
			32'd712:
				output_byte = 8'd0;
			32'd713:
				output_byte = 8'd0;
			32'd714:
				output_byte = 8'd0;
			32'd715:
				output_byte = 8'd8;
			32'd716:
				output_byte = 8'd3;
			32'd717:
				output_byte = 8'd0;
			32'd718:
				output_byte = 8'd0;
			32'd719:
				output_byte = 8'd0;
			32'd720:
				output_byte = 8'd1;
			32'd721:
				output_byte = 8'd0;
			32'd722:
				output_byte = 8'd0;
			32'd723:
				output_byte = 8'd0;
			32'd724:
				output_byte = 8'd10;
			32'd725:
				output_byte = 8'd235;
			32'd726:
				output_byte = 8'd2;
			32'd727:
				output_byte = 8'd0;
			32'd728:
				output_byte = 8'd0;
			32'd729:
				output_byte = 8'd0;
			32'd730:
				output_byte = 8'd0;
			32'd731:
				output_byte = 8'd0;
			32'd732:
				output_byte = 8'd0;
			32'd733:
				output_byte = 8'd9;
			32'd734:
				output_byte = 8'd235;
			32'd735:
				output_byte = 8'd2;
			32'd736:
				output_byte = 8'd0;
			32'd737:
				output_byte = 8'd0;
			32'd738:
				output_byte = 8'd0;
			32'd739:
				output_byte = 8'd0;
			32'd740:
				output_byte = 8'd0;
			32'd741:
				output_byte = 8'd0;
			32'd742:
				output_byte = 8'd20;
			32'd743:
				output_byte = 8'd0;
			32'd744:
				output_byte = 8'd0;
			32'd745:
				output_byte = 8'd0;
			32'd746:
				output_byte = 8'd0;
			32'd747:
				output_byte = 8'd1;
			32'd748:
				output_byte = 8'd0;
			32'd749:
				output_byte = 8'd0;
			32'd750:
				output_byte = 8'd0;
			32'd751:
				output_byte = 8'd1;
			32'd752:
				output_byte = 8'd24;
			32'd753:
				output_byte = 8'd0;
			32'd754:
				output_byte = 8'd0;
			32'd755:
				output_byte = 8'd0;
			32'd756:
				output_byte = 8'd2;
			32'd757:
				output_byte = 8'd0;
			32'd758:
				output_byte = 8'd0;
			32'd759:
				output_byte = 8'd0;
			32'd760:
				output_byte = 8'd3;
			32'd761:
				output_byte = 8'd1;
			32'd762:
				output_byte = 8'd0;
			32'd763:
				output_byte = 8'd0;
			32'd764:
				output_byte = 8'd0;
			32'd765:
				output_byte = 8'd2;
			32'd766:
				output_byte = 8'd0;
			32'd767:
				output_byte = 8'd0;
			32'd768:
				output_byte = 8'd0;
			32'd769:
				output_byte = 8'd20;
			32'd770:
				output_byte = 8'd1;
			32'd771:
				output_byte = 8'd0;
			32'd772:
				output_byte = 8'd0;
			32'd773:
				output_byte = 8'd0;
			32'd774:
				output_byte = 8'd2;
			32'd775:
				output_byte = 8'd0;
			32'd776:
				output_byte = 8'd0;
			32'd777:
				output_byte = 8'd0;
			32'd778:
				output_byte = 8'd3;
			32'd779:
				output_byte = 8'd1;
			32'd780:
				output_byte = 8'd0;
			32'd781:
				output_byte = 8'd0;
			32'd782:
				output_byte = 8'd0;
			32'd783:
				output_byte = 8'd2;
			32'd784:
				output_byte = 8'd0;
			32'd785:
				output_byte = 8'd0;
			32'd786:
				output_byte = 8'd0;
			32'd787:
				output_byte = 8'd2;
			32'd788:
				output_byte = 8'd1;
			32'd789:
				output_byte = 8'd0;
			32'd790:
				output_byte = 8'd0;
			32'd791:
				output_byte = 8'd0;
			32'd792:
				output_byte = 8'd24;
			32'd793:
				output_byte = 8'd0;
			32'd794:
				output_byte = 8'd0;
			32'd795:
				output_byte = 8'd0;
			32'd796:
				output_byte = 8'd8;
			32'd797:
				output_byte = 8'd1;
			32'd798:
				output_byte = 8'd0;
			32'd799:
				output_byte = 8'd0;
			32'd800:
				output_byte = 8'd0;
			32'd801:
				output_byte = 8'd1;
			32'd802:
				output_byte = 8'd0;
			32'd803:
				output_byte = 8'd0;
			32'd804:
				output_byte = 8'd0;
			32'd805:
				output_byte = 8'd10;
			32'd806:
				output_byte = 8'd32;
			32'd807:
				output_byte = 8'd1;
			32'd808:
				output_byte = 8'd0;
			32'd809:
				output_byte = 8'd0;
			32'd810:
				output_byte = 8'd0;
			32'd811:
				output_byte = 8'd0;
			32'd812:
				output_byte = 8'd0;
			32'd813:
				output_byte = 8'd0;
			32'd814:
				output_byte = 8'd20;
			32'd815:
				output_byte = 8'd0;
			32'd816:
				output_byte = 8'd0;
			32'd817:
				output_byte = 8'd0;
			32'd818:
				output_byte = 8'd0;
			32'd819:
				output_byte = 8'd1;
			32'd820:
				output_byte = 8'd0;
			32'd821:
				output_byte = 8'd0;
			32'd822:
				output_byte = 8'd0;
			32'd823:
				output_byte = 8'd1;
			32'd824:
				output_byte = 8'd32;
			32'd825:
				output_byte = 8'd0;
			32'd826:
				output_byte = 8'd0;
			32'd827:
				output_byte = 8'd0;
			32'd828:
				output_byte = 8'd2;
			32'd829:
				output_byte = 8'd0;
			32'd830:
				output_byte = 8'd0;
			32'd831:
				output_byte = 8'd0;
			32'd832:
				output_byte = 8'd3;
			32'd833:
				output_byte = 8'd1;
			32'd834:
				output_byte = 8'd0;
			32'd835:
				output_byte = 8'd0;
			32'd836:
				output_byte = 8'd0;
			32'd837:
				output_byte = 8'd2;
			32'd838:
				output_byte = 8'd0;
			32'd839:
				output_byte = 8'd0;
			32'd840:
				output_byte = 8'd0;
			32'd841:
				output_byte = 8'd7;
			32'd842:
				output_byte = 8'd1;
			32'd843:
				output_byte = 8'd0;
			32'd844:
				output_byte = 8'd0;
			32'd845:
				output_byte = 8'd0;
			32'd846:
				output_byte = 8'd3;
			32'd847:
				output_byte = 8'd0;
			32'd848:
				output_byte = 8'd0;
			32'd849:
				output_byte = 8'd0;
			32'd850:
				output_byte = 8'd20;
			32'd851:
				output_byte = 8'd0;
			32'd852:
				output_byte = 8'd0;
			32'd853:
				output_byte = 8'd0;
			32'd854:
				output_byte = 8'd0;
			32'd855:
				output_byte = 8'd1;
			32'd856:
				output_byte = 8'd0;
			32'd857:
				output_byte = 8'd0;
			32'd858:
				output_byte = 8'd0;
			32'd859:
				output_byte = 8'd20;
			32'd860:
				output_byte = 8'd1;
			32'd861:
				output_byte = 8'd0;
			32'd862:
				output_byte = 8'd0;
			32'd863:
				output_byte = 8'd0;
			32'd864:
				output_byte = 8'd2;
			32'd865:
				output_byte = 8'd0;
			32'd866:
				output_byte = 8'd0;
			32'd867:
				output_byte = 8'd0;
			32'd868:
				output_byte = 8'd3;
			32'd869:
				output_byte = 8'd1;
			32'd870:
				output_byte = 8'd0;
			32'd871:
				output_byte = 8'd0;
			32'd872:
				output_byte = 8'd0;
			32'd873:
				output_byte = 8'd2;
			32'd874:
				output_byte = 8'd0;
			32'd875:
				output_byte = 8'd0;
			32'd876:
				output_byte = 8'd0;
			32'd877:
				output_byte = 8'd8;
			32'd878:
				output_byte = 8'd3;
			32'd879:
				output_byte = 8'd0;
			32'd880:
				output_byte = 8'd0;
			32'd881:
				output_byte = 8'd0;
			32'd882:
				output_byte = 8'd1;
			32'd883:
				output_byte = 8'd0;
			32'd884:
				output_byte = 8'd0;
			32'd885:
				output_byte = 8'd0;
			32'd886:
				output_byte = 8'd9;
			32'd887:
				output_byte = 8'd201;
			32'd888:
				output_byte = 8'd6;
			32'd889:
				output_byte = 8'd0;
			32'd890:
				output_byte = 8'd0;
			32'd891:
				output_byte = 8'd0;
			32'd892:
				output_byte = 8'd0;
			32'd893:
				output_byte = 8'd0;
			32'd894:
				output_byte = 8'd0;
			32'd895:
				output_byte = 8'd11;
			32'd896:
				output_byte = 8'd201;
			32'd897:
				output_byte = 8'd6;
			32'd898:
				output_byte = 8'd0;
			32'd899:
				output_byte = 8'd0;
			32'd900:
				output_byte = 8'd0;
			32'd901:
				output_byte = 8'd0;
			32'd902:
				output_byte = 8'd0;
			32'd903:
				output_byte = 8'd0;
			32'd904:
				output_byte = 8'd20;
			32'd905:
				output_byte = 8'd0;
			32'd906:
				output_byte = 8'd0;
			32'd907:
				output_byte = 8'd0;
			32'd908:
				output_byte = 8'd0;
			32'd909:
				output_byte = 8'd1;
			32'd910:
				output_byte = 8'd0;
			32'd911:
				output_byte = 8'd0;
			32'd912:
				output_byte = 8'd0;
			32'd913:
				output_byte = 8'd2;
			32'd914:
				output_byte = 8'd1;
			32'd915:
				output_byte = 8'd0;
			32'd916:
				output_byte = 8'd0;
			32'd917:
				output_byte = 8'd0;
			32'd918:
				output_byte = 8'd36;
			32'd919:
				output_byte = 8'd0;
			32'd920:
				output_byte = 8'd0;
			32'd921:
				output_byte = 8'd0;
			32'd922:
				output_byte = 8'd20;
			32'd923:
				output_byte = 8'd0;
			32'd924:
				output_byte = 8'd0;
			32'd925:
				output_byte = 8'd0;
			32'd926:
				output_byte = 8'd0;
			32'd927:
				output_byte = 8'd1;
			32'd928:
				output_byte = 8'd0;
			32'd929:
				output_byte = 8'd0;
			32'd930:
				output_byte = 8'd0;
			32'd931:
				output_byte = 8'd2;
			32'd932:
				output_byte = 8'd1;
			32'd933:
				output_byte = 8'd0;
			32'd934:
				output_byte = 8'd0;
			32'd935:
				output_byte = 8'd0;
			32'd936:
				output_byte = 8'd40;
			32'd937:
				output_byte = 8'd0;
			32'd938:
				output_byte = 8'd0;
			32'd939:
				output_byte = 8'd0;
			32'd940:
				output_byte = 8'd20;
			32'd941:
				output_byte = 8'd0;
			32'd942:
				output_byte = 8'd0;
			32'd943:
				output_byte = 8'd0;
			32'd944:
				output_byte = 8'd0;
			32'd945:
				output_byte = 8'd1;
			32'd946:
				output_byte = 8'd0;
			32'd947:
				output_byte = 8'd0;
			32'd948:
				output_byte = 8'd0;
			32'd949:
				output_byte = 8'd1;
			32'd950:
				output_byte = 8'd16;
			32'd951:
				output_byte = 8'd0;
			32'd952:
				output_byte = 8'd0;
			32'd953:
				output_byte = 8'd0;
			32'd954:
				output_byte = 8'd2;
			32'd955:
				output_byte = 8'd0;
			32'd956:
				output_byte = 8'd0;
			32'd957:
				output_byte = 8'd0;
			32'd958:
				output_byte = 8'd3;
			32'd959:
				output_byte = 8'd1;
			32'd960:
				output_byte = 8'd0;
			32'd961:
				output_byte = 8'd0;
			32'd962:
				output_byte = 8'd0;
			32'd963:
				output_byte = 8'd2;
			32'd964:
				output_byte = 8'd0;
			32'd965:
				output_byte = 8'd0;
			32'd966:
				output_byte = 8'd0;
			32'd967:
				output_byte = 8'd2;
			32'd968:
				output_byte = 8'd1;
			32'd969:
				output_byte = 8'd0;
			32'd970:
				output_byte = 8'd0;
			32'd971:
				output_byte = 8'd0;
			32'd972:
				output_byte = 8'd40;
			32'd973:
				output_byte = 8'd0;
			32'd974:
				output_byte = 8'd0;
			32'd975:
				output_byte = 8'd0;
			32'd976:
				output_byte = 8'd20;
			32'd977:
				output_byte = 8'd0;
			32'd978:
				output_byte = 8'd0;
			32'd979:
				output_byte = 8'd0;
			32'd980:
				output_byte = 8'd0;
			32'd981:
				output_byte = 8'd1;
			32'd982:
				output_byte = 8'd0;
			32'd983:
				output_byte = 8'd0;
			32'd984:
				output_byte = 8'd0;
			32'd985:
				output_byte = 8'd1;
			32'd986:
				output_byte = 8'd40;
			32'd987:
				output_byte = 8'd0;
			32'd988:
				output_byte = 8'd0;
			32'd989:
				output_byte = 8'd0;
			32'd990:
				output_byte = 8'd2;
			32'd991:
				output_byte = 8'd0;
			32'd992:
				output_byte = 8'd0;
			32'd993:
				output_byte = 8'd0;
			32'd994:
				output_byte = 8'd3;
			32'd995:
				output_byte = 8'd1;
			32'd996:
				output_byte = 8'd0;
			32'd997:
				output_byte = 8'd0;
			32'd998:
				output_byte = 8'd0;
			32'd999:
				output_byte = 8'd2;
			32'd1000:
				output_byte = 8'd0;
			32'd1001:
				output_byte = 8'd0;
			32'd1002:
				output_byte = 8'd0;
			32'd1003:
				output_byte = 8'd7;
			32'd1004:
				output_byte = 8'd1;
			32'd1005:
				output_byte = 8'd0;
			32'd1006:
				output_byte = 8'd0;
			32'd1007:
				output_byte = 8'd0;
			32'd1008:
				output_byte = 8'd3;
			32'd1009:
				output_byte = 8'd0;
			32'd1010:
				output_byte = 8'd0;
			32'd1011:
				output_byte = 8'd0;
			32'd1012:
				output_byte = 8'd20;
			32'd1013:
				output_byte = 8'd0;
			32'd1014:
				output_byte = 8'd0;
			32'd1015:
				output_byte = 8'd0;
			32'd1016:
				output_byte = 8'd0;
			32'd1017:
				output_byte = 8'd1;
			32'd1018:
				output_byte = 8'd0;
			32'd1019:
				output_byte = 8'd0;
			32'd1020:
				output_byte = 8'd0;
			32'd1021:
				output_byte = 8'd20;
			32'd1022:
				output_byte = 8'd0;
			32'd1023:
				output_byte = 8'd0;
			32'd1024:
				output_byte = 8'd0;
			32'd1025:
				output_byte = 8'd0;
			32'd1026:
				output_byte = 8'd2;
			32'd1027:
				output_byte = 8'd0;
			32'd1028:
				output_byte = 8'd0;
			32'd1029:
				output_byte = 8'd0;
			32'd1030:
				output_byte = 8'd3;
			32'd1031:
				output_byte = 8'd1;
			32'd1032:
				output_byte = 8'd0;
			32'd1033:
				output_byte = 8'd0;
			32'd1034:
				output_byte = 8'd0;
			32'd1035:
				output_byte = 8'd2;
			32'd1036:
				output_byte = 8'd0;
			32'd1037:
				output_byte = 8'd0;
			32'd1038:
				output_byte = 8'd0;
			32'd1039:
				output_byte = 8'd8;
			32'd1040:
				output_byte = 8'd3;
			32'd1041:
				output_byte = 8'd0;
			32'd1042:
				output_byte = 8'd0;
			32'd1043:
				output_byte = 8'd0;
			32'd1044:
				output_byte = 8'd1;
			32'd1045:
				output_byte = 8'd0;
			32'd1046:
				output_byte = 8'd0;
			32'd1047:
				output_byte = 8'd0;
			32'd1048:
				output_byte = 8'd10;
			32'd1049:
				output_byte = 8'd119;
			32'd1050:
				output_byte = 8'd4;
			32'd1051:
				output_byte = 8'd0;
			32'd1052:
				output_byte = 8'd0;
			32'd1053:
				output_byte = 8'd0;
			32'd1054:
				output_byte = 8'd0;
			32'd1055:
				output_byte = 8'd0;
			32'd1056:
				output_byte = 8'd0;
			32'd1057:
				output_byte = 8'd9;
			32'd1058:
				output_byte = 8'd119;
			32'd1059:
				output_byte = 8'd4;
			32'd1060:
				output_byte = 8'd0;
			32'd1061:
				output_byte = 8'd0;
			32'd1062:
				output_byte = 8'd0;
			32'd1063:
				output_byte = 8'd0;
			32'd1064:
				output_byte = 8'd0;
			32'd1065:
				output_byte = 8'd0;
			32'd1066:
				output_byte = 8'd20;
			32'd1067:
				output_byte = 8'd0;
			32'd1068:
				output_byte = 8'd0;
			32'd1069:
				output_byte = 8'd0;
			32'd1070:
				output_byte = 8'd0;
			32'd1071:
				output_byte = 8'd1;
			32'd1072:
				output_byte = 8'd0;
			32'd1073:
				output_byte = 8'd0;
			32'd1074:
				output_byte = 8'd0;
			32'd1075:
				output_byte = 8'd1;
			32'd1076:
				output_byte = 8'd40;
			32'd1077:
				output_byte = 8'd0;
			32'd1078:
				output_byte = 8'd0;
			32'd1079:
				output_byte = 8'd0;
			32'd1080:
				output_byte = 8'd2;
			32'd1081:
				output_byte = 8'd0;
			32'd1082:
				output_byte = 8'd0;
			32'd1083:
				output_byte = 8'd0;
			32'd1084:
				output_byte = 8'd3;
			32'd1085:
				output_byte = 8'd1;
			32'd1086:
				output_byte = 8'd0;
			32'd1087:
				output_byte = 8'd0;
			32'd1088:
				output_byte = 8'd0;
			32'd1089:
				output_byte = 8'd2;
			32'd1090:
				output_byte = 8'd0;
			32'd1091:
				output_byte = 8'd0;
			32'd1092:
				output_byte = 8'd0;
			32'd1093:
				output_byte = 8'd20;
			32'd1094:
				output_byte = 8'd10;
			32'd1095:
				output_byte = 8'd0;
			32'd1096:
				output_byte = 8'd0;
			32'd1097:
				output_byte = 8'd0;
			32'd1098:
				output_byte = 8'd2;
			32'd1099:
				output_byte = 8'd0;
			32'd1100:
				output_byte = 8'd0;
			32'd1101:
				output_byte = 8'd0;
			32'd1102:
				output_byte = 8'd22;
			32'd1103:
				output_byte = 8'd1;
			32'd1104:
				output_byte = 8'd0;
			32'd1105:
				output_byte = 8'd0;
			32'd1106:
				output_byte = 8'd0;
			32'd1107:
				output_byte = 8'd2;
			32'd1108:
				output_byte = 8'd0;
			32'd1109:
				output_byte = 8'd0;
			32'd1110:
				output_byte = 8'd0;
			32'd1111:
				output_byte = 8'd2;
			32'd1112:
				output_byte = 8'd1;
			32'd1113:
				output_byte = 8'd0;
			32'd1114:
				output_byte = 8'd0;
			32'd1115:
				output_byte = 8'd0;
			32'd1116:
				output_byte = 8'd40;
			32'd1117:
				output_byte = 8'd0;
			32'd1118:
				output_byte = 8'd0;
			32'd1119:
				output_byte = 8'd0;
			32'd1120:
				output_byte = 8'd20;
			32'd1121:
				output_byte = 8'd0;
			32'd1122:
				output_byte = 8'd0;
			32'd1123:
				output_byte = 8'd0;
			32'd1124:
				output_byte = 8'd0;
			32'd1125:
				output_byte = 8'd1;
			32'd1126:
				output_byte = 8'd0;
			32'd1127:
				output_byte = 8'd0;
			32'd1128:
				output_byte = 8'd0;
			32'd1129:
				output_byte = 8'd1;
			32'd1130:
				output_byte = 8'd36;
			32'd1131:
				output_byte = 8'd0;
			32'd1132:
				output_byte = 8'd0;
			32'd1133:
				output_byte = 8'd0;
			32'd1134:
				output_byte = 8'd2;
			32'd1135:
				output_byte = 8'd0;
			32'd1136:
				output_byte = 8'd0;
			32'd1137:
				output_byte = 8'd0;
			32'd1138:
				output_byte = 8'd3;
			32'd1139:
				output_byte = 8'd1;
			32'd1140:
				output_byte = 8'd0;
			32'd1141:
				output_byte = 8'd0;
			32'd1142:
				output_byte = 8'd0;
			32'd1143:
				output_byte = 8'd2;
			32'd1144:
				output_byte = 8'd0;
			32'd1145:
				output_byte = 8'd0;
			32'd1146:
				output_byte = 8'd0;
			32'd1147:
				output_byte = 8'd20;
			32'd1148:
				output_byte = 8'd1;
			32'd1149:
				output_byte = 8'd0;
			32'd1150:
				output_byte = 8'd0;
			32'd1151:
				output_byte = 8'd0;
			32'd1152:
				output_byte = 8'd2;
			32'd1153:
				output_byte = 8'd0;
			32'd1154:
				output_byte = 8'd0;
			32'd1155:
				output_byte = 8'd0;
			32'd1156:
				output_byte = 8'd3;
			32'd1157:
				output_byte = 8'd1;
			32'd1158:
				output_byte = 8'd0;
			32'd1159:
				output_byte = 8'd0;
			32'd1160:
				output_byte = 8'd0;
			32'd1161:
				output_byte = 8'd2;
			32'd1162:
				output_byte = 8'd0;
			32'd1163:
				output_byte = 8'd0;
			32'd1164:
				output_byte = 8'd0;
			32'd1165:
				output_byte = 8'd2;
			32'd1166:
				output_byte = 8'd1;
			32'd1167:
				output_byte = 8'd0;
			32'd1168:
				output_byte = 8'd0;
			32'd1169:
				output_byte = 8'd0;
			32'd1170:
				output_byte = 8'd36;
			32'd1171:
				output_byte = 8'd0;
			32'd1172:
				output_byte = 8'd0;
			32'd1173:
				output_byte = 8'd0;
			32'd1174:
				output_byte = 8'd8;
			32'd1175:
				output_byte = 8'd1;
			32'd1176:
				output_byte = 8'd0;
			32'd1177:
				output_byte = 8'd0;
			32'd1178:
				output_byte = 8'd0;
			32'd1179:
				output_byte = 8'd1;
			32'd1180:
				output_byte = 8'd0;
			32'd1181:
				output_byte = 8'd0;
			32'd1182:
				output_byte = 8'd0;
			32'd1183:
				output_byte = 8'd10;
			32'd1184:
				output_byte = 8'd159;
			32'd1185:
				output_byte = 8'd3;
			32'd1186:
				output_byte = 8'd0;
			32'd1187:
				output_byte = 8'd0;
			32'd1188:
				output_byte = 8'd0;
			32'd1189:
				output_byte = 8'd0;
			32'd1190:
				output_byte = 8'd0;
			32'd1191:
				output_byte = 8'd0;
			32'd1192:
				output_byte = 8'd20;
			32'd1193:
				output_byte = 8'd0;
			32'd1194:
				output_byte = 8'd0;
			32'd1195:
				output_byte = 8'd0;
			32'd1196:
				output_byte = 8'd0;
			32'd1197:
				output_byte = 8'd1;
			32'd1198:
				output_byte = 8'd0;
			32'd1199:
				output_byte = 8'd0;
			32'd1200:
				output_byte = 8'd0;
			32'd1201:
				output_byte = 8'd1;
			32'd1202:
				output_byte = 8'd16;
			32'd1203:
				output_byte = 8'd0;
			32'd1204:
				output_byte = 8'd0;
			32'd1205:
				output_byte = 8'd0;
			32'd1206:
				output_byte = 8'd2;
			32'd1207:
				output_byte = 8'd0;
			32'd1208:
				output_byte = 8'd0;
			32'd1209:
				output_byte = 8'd0;
			32'd1210:
				output_byte = 8'd3;
			32'd1211:
				output_byte = 8'd1;
			32'd1212:
				output_byte = 8'd0;
			32'd1213:
				output_byte = 8'd0;
			32'd1214:
				output_byte = 8'd0;
			32'd1215:
				output_byte = 8'd2;
			32'd1216:
				output_byte = 8'd0;
			32'd1217:
				output_byte = 8'd0;
			32'd1218:
				output_byte = 8'd0;
			32'd1219:
				output_byte = 8'd2;
			32'd1220:
				output_byte = 8'd1;
			32'd1221:
				output_byte = 8'd0;
			32'd1222:
				output_byte = 8'd0;
			32'd1223:
				output_byte = 8'd0;
			32'd1224:
				output_byte = 8'd40;
			32'd1225:
				output_byte = 8'd0;
			32'd1226:
				output_byte = 8'd0;
			32'd1227:
				output_byte = 8'd0;
			32'd1228:
				output_byte = 8'd20;
			32'd1229:
				output_byte = 8'd0;
			32'd1230:
				output_byte = 8'd0;
			32'd1231:
				output_byte = 8'd0;
			32'd1232:
				output_byte = 8'd0;
			32'd1233:
				output_byte = 8'd1;
			32'd1234:
				output_byte = 8'd0;
			32'd1235:
				output_byte = 8'd0;
			32'd1236:
				output_byte = 8'd0;
			32'd1237:
				output_byte = 8'd1;
			32'd1238:
				output_byte = 8'd40;
			32'd1239:
				output_byte = 8'd0;
			32'd1240:
				output_byte = 8'd0;
			32'd1241:
				output_byte = 8'd0;
			32'd1242:
				output_byte = 8'd2;
			32'd1243:
				output_byte = 8'd0;
			32'd1244:
				output_byte = 8'd0;
			32'd1245:
				output_byte = 8'd0;
			32'd1246:
				output_byte = 8'd3;
			32'd1247:
				output_byte = 8'd1;
			32'd1248:
				output_byte = 8'd0;
			32'd1249:
				output_byte = 8'd0;
			32'd1250:
				output_byte = 8'd0;
			32'd1251:
				output_byte = 8'd2;
			32'd1252:
				output_byte = 8'd0;
			32'd1253:
				output_byte = 8'd0;
			32'd1254:
				output_byte = 8'd0;
			32'd1255:
				output_byte = 8'd7;
			32'd1256:
				output_byte = 8'd1;
			32'd1257:
				output_byte = 8'd0;
			32'd1258:
				output_byte = 8'd0;
			32'd1259:
				output_byte = 8'd0;
			32'd1260:
				output_byte = 8'd3;
			32'd1261:
				output_byte = 8'd0;
			32'd1262:
				output_byte = 8'd0;
			32'd1263:
				output_byte = 8'd0;
			32'd1264:
				output_byte = 8'd20;
			32'd1265:
				output_byte = 8'd0;
			32'd1266:
				output_byte = 8'd0;
			32'd1267:
				output_byte = 8'd0;
			32'd1268:
				output_byte = 8'd0;
			32'd1269:
				output_byte = 8'd1;
			32'd1270:
				output_byte = 8'd0;
			32'd1271:
				output_byte = 8'd0;
			32'd1272:
				output_byte = 8'd0;
			32'd1273:
				output_byte = 8'd20;
			32'd1274:
				output_byte = 8'd0;
			32'd1275:
				output_byte = 8'd0;
			32'd1276:
				output_byte = 8'd0;
			32'd1277:
				output_byte = 8'd0;
			32'd1278:
				output_byte = 8'd2;
			32'd1279:
				output_byte = 8'd0;
			32'd1280:
				output_byte = 8'd0;
			32'd1281:
				output_byte = 8'd0;
			32'd1282:
				output_byte = 8'd3;
			32'd1283:
				output_byte = 8'd1;
			32'd1284:
				output_byte = 8'd0;
			32'd1285:
				output_byte = 8'd0;
			32'd1286:
				output_byte = 8'd0;
			32'd1287:
				output_byte = 8'd2;
			32'd1288:
				output_byte = 8'd0;
			32'd1289:
				output_byte = 8'd0;
			32'd1290:
				output_byte = 8'd0;
			32'd1291:
				output_byte = 8'd8;
			32'd1292:
				output_byte = 8'd3;
			32'd1293:
				output_byte = 8'd0;
			32'd1294:
				output_byte = 8'd0;
			32'd1295:
				output_byte = 8'd0;
			32'd1296:
				output_byte = 8'd1;
			32'd1297:
				output_byte = 8'd0;
			32'd1298:
				output_byte = 8'd0;
			32'd1299:
				output_byte = 8'd0;
			32'd1300:
				output_byte = 8'd10;
			32'd1301:
				output_byte = 8'd147;
			32'd1302:
				output_byte = 8'd6;
			32'd1303:
				output_byte = 8'd0;
			32'd1304:
				output_byte = 8'd0;
			32'd1305:
				output_byte = 8'd0;
			32'd1306:
				output_byte = 8'd0;
			32'd1307:
				output_byte = 8'd0;
			32'd1308:
				output_byte = 8'd0;
			32'd1309:
				output_byte = 8'd9;
			32'd1310:
				output_byte = 8'd147;
			32'd1311:
				output_byte = 8'd6;
			32'd1312:
				output_byte = 8'd0;
			32'd1313:
				output_byte = 8'd0;
			32'd1314:
				output_byte = 8'd0;
			32'd1315:
				output_byte = 8'd0;
			32'd1316:
				output_byte = 8'd0;
			32'd1317:
				output_byte = 8'd0;
			32'd1318:
				output_byte = 8'd20;
			32'd1319:
				output_byte = 8'd0;
			32'd1320:
				output_byte = 8'd0;
			32'd1321:
				output_byte = 8'd0;
			32'd1322:
				output_byte = 8'd0;
			32'd1323:
				output_byte = 8'd1;
			32'd1324:
				output_byte = 8'd0;
			32'd1325:
				output_byte = 8'd0;
			32'd1326:
				output_byte = 8'd0;
			32'd1327:
				output_byte = 8'd2;
			32'd1328:
				output_byte = 8'd1;
			32'd1329:
				output_byte = 8'd0;
			32'd1330:
				output_byte = 8'd0;
			32'd1331:
				output_byte = 8'd0;
			32'd1332:
				output_byte = 8'd44;
			32'd1333:
				output_byte = 8'd0;
			32'd1334:
				output_byte = 8'd0;
			32'd1335:
				output_byte = 8'd0;
			32'd1336:
				output_byte = 8'd20;
			32'd1337:
				output_byte = 8'd0;
			32'd1338:
				output_byte = 8'd0;
			32'd1339:
				output_byte = 8'd0;
			32'd1340:
				output_byte = 8'd0;
			32'd1341:
				output_byte = 8'd1;
			32'd1342:
				output_byte = 8'd0;
			32'd1343:
				output_byte = 8'd0;
			32'd1344:
				output_byte = 8'd0;
			32'd1345:
				output_byte = 8'd1;
			32'd1346:
				output_byte = 8'd40;
			32'd1347:
				output_byte = 8'd0;
			32'd1348:
				output_byte = 8'd0;
			32'd1349:
				output_byte = 8'd0;
			32'd1350:
				output_byte = 8'd2;
			32'd1351:
				output_byte = 8'd0;
			32'd1352:
				output_byte = 8'd0;
			32'd1353:
				output_byte = 8'd0;
			32'd1354:
				output_byte = 8'd3;
			32'd1355:
				output_byte = 8'd1;
			32'd1356:
				output_byte = 8'd0;
			32'd1357:
				output_byte = 8'd0;
			32'd1358:
				output_byte = 8'd0;
			32'd1359:
				output_byte = 8'd2;
			32'd1360:
				output_byte = 8'd0;
			32'd1361:
				output_byte = 8'd0;
			32'd1362:
				output_byte = 8'd0;
			32'd1363:
				output_byte = 8'd20;
			32'd1364:
				output_byte = 8'd10;
			32'd1365:
				output_byte = 8'd0;
			32'd1366:
				output_byte = 8'd0;
			32'd1367:
				output_byte = 8'd0;
			32'd1368:
				output_byte = 8'd2;
			32'd1369:
				output_byte = 8'd0;
			32'd1370:
				output_byte = 8'd0;
			32'd1371:
				output_byte = 8'd0;
			32'd1372:
				output_byte = 8'd22;
			32'd1373:
				output_byte = 8'd1;
			32'd1374:
				output_byte = 8'd0;
			32'd1375:
				output_byte = 8'd0;
			32'd1376:
				output_byte = 8'd0;
			32'd1377:
				output_byte = 8'd2;
			32'd1378:
				output_byte = 8'd0;
			32'd1379:
				output_byte = 8'd0;
			32'd1380:
				output_byte = 8'd0;
			32'd1381:
				output_byte = 8'd7;
			32'd1382:
				output_byte = 8'd2;
			32'd1383:
				output_byte = 8'd0;
			32'd1384:
				output_byte = 8'd0;
			32'd1385:
				output_byte = 8'd0;
			32'd1386:
				output_byte = 8'd1;
			32'd1387:
				output_byte = 8'd0;
			32'd1388:
				output_byte = 8'd0;
			32'd1389:
				output_byte = 8'd0;
			32'd1390:
				output_byte = 8'd2;
			32'd1391:
				output_byte = 8'd1;
			32'd1392:
				output_byte = 8'd0;
			32'd1393:
				output_byte = 8'd0;
			32'd1394:
				output_byte = 8'd0;
			32'd1395:
				output_byte = 8'd44;
			32'd1396:
				output_byte = 8'd0;
			32'd1397:
				output_byte = 8'd0;
			32'd1398:
				output_byte = 8'd0;
			32'd1399:
				output_byte = 8'd20;
			32'd1400:
				output_byte = 8'd0;
			32'd1401:
				output_byte = 8'd0;
			32'd1402:
				output_byte = 8'd0;
			32'd1403:
				output_byte = 8'd0;
			32'd1404:
				output_byte = 8'd1;
			32'd1405:
				output_byte = 8'd0;
			32'd1406:
				output_byte = 8'd0;
			32'd1407:
				output_byte = 8'd0;
			32'd1408:
				output_byte = 8'd1;
			32'd1409:
				output_byte = 8'd12;
			32'd1410:
				output_byte = 8'd0;
			32'd1411:
				output_byte = 8'd0;
			32'd1412:
				output_byte = 8'd0;
			32'd1413:
				output_byte = 8'd2;
			32'd1414:
				output_byte = 8'd0;
			32'd1415:
				output_byte = 8'd0;
			32'd1416:
				output_byte = 8'd0;
			32'd1417:
				output_byte = 8'd3;
			32'd1418:
				output_byte = 8'd1;
			32'd1419:
				output_byte = 8'd0;
			32'd1420:
				output_byte = 8'd0;
			32'd1421:
				output_byte = 8'd0;
			32'd1422:
				output_byte = 8'd2;
			32'd1423:
				output_byte = 8'd0;
			32'd1424:
				output_byte = 8'd0;
			32'd1425:
				output_byte = 8'd0;
			32'd1426:
				output_byte = 8'd1;
			32'd1427:
				output_byte = 8'd20;
			32'd1428:
				output_byte = 8'd0;
			32'd1429:
				output_byte = 8'd0;
			32'd1430:
				output_byte = 8'd0;
			32'd1431:
				output_byte = 8'd2;
			32'd1432:
				output_byte = 8'd0;
			32'd1433:
				output_byte = 8'd0;
			32'd1434:
				output_byte = 8'd0;
			32'd1435:
				output_byte = 8'd21;
			32'd1436:
				output_byte = 8'd1;
			32'd1437:
				output_byte = 8'd0;
			32'd1438:
				output_byte = 8'd0;
			32'd1439:
				output_byte = 8'd0;
			32'd1440:
				output_byte = 8'd2;
			32'd1441:
				output_byte = 8'd0;
			32'd1442:
				output_byte = 8'd0;
			32'd1443:
				output_byte = 8'd0;
			32'd1444:
				output_byte = 8'd2;
			32'd1445:
				output_byte = 8'd1;
			32'd1446:
				output_byte = 8'd0;
			32'd1447:
				output_byte = 8'd0;
			32'd1448:
				output_byte = 8'd0;
			32'd1449:
				output_byte = 8'd0;
			32'd1450:
				output_byte = 8'd0;
			32'd1451:
				output_byte = 8'd0;
			32'd1452:
				output_byte = 8'd0;
			32'd1453:
				output_byte = 8'd20;
			32'd1454:
				output_byte = 8'd0;
			32'd1455:
				output_byte = 8'd0;
			32'd1456:
				output_byte = 8'd0;
			32'd1457:
				output_byte = 8'd0;
			32'd1458:
				output_byte = 8'd1;
			32'd1459:
				output_byte = 8'd0;
			32'd1460:
				output_byte = 8'd0;
			32'd1461:
				output_byte = 8'd0;
			32'd1462:
				output_byte = 8'd1;
			32'd1463:
				output_byte = 8'd0;
			32'd1464:
				output_byte = 8'd0;
			32'd1465:
				output_byte = 8'd0;
			32'd1466:
				output_byte = 8'd0;
			32'd1467:
				output_byte = 8'd2;
			32'd1468:
				output_byte = 8'd0;
			32'd1469:
				output_byte = 8'd0;
			32'd1470:
				output_byte = 8'd0;
			32'd1471:
				output_byte = 8'd3;
			32'd1472:
				output_byte = 8'd1;
			32'd1473:
				output_byte = 8'd0;
			32'd1474:
				output_byte = 8'd0;
			32'd1475:
				output_byte = 8'd0;
			32'd1476:
				output_byte = 8'd2;
			32'd1477:
				output_byte = 8'd0;
			32'd1478:
				output_byte = 8'd0;
			32'd1479:
				output_byte = 8'd0;
			32'd1480:
				output_byte = 8'd1;
			32'd1481:
				output_byte = 8'd36;
			32'd1482:
				output_byte = 8'd0;
			32'd1483:
				output_byte = 8'd0;
			32'd1484:
				output_byte = 8'd0;
			32'd1485:
				output_byte = 8'd2;
			32'd1486:
				output_byte = 8'd0;
			32'd1487:
				output_byte = 8'd0;
			32'd1488:
				output_byte = 8'd0;
			32'd1489:
				output_byte = 8'd3;
			32'd1490:
				output_byte = 8'd1;
			32'd1491:
				output_byte = 8'd0;
			32'd1492:
				output_byte = 8'd0;
			32'd1493:
				output_byte = 8'd0;
			32'd1494:
				output_byte = 8'd2;
			32'd1495:
				output_byte = 8'd0;
			32'd1496:
				output_byte = 8'd0;
			32'd1497:
				output_byte = 8'd0;
			32'd1498:
				output_byte = 8'd20;
			32'd1499:
				output_byte = 8'd1;
			32'd1500:
				output_byte = 8'd0;
			32'd1501:
				output_byte = 8'd0;
			32'd1502:
				output_byte = 8'd0;
			32'd1503:
				output_byte = 8'd2;
			32'd1504:
				output_byte = 8'd0;
			32'd1505:
				output_byte = 8'd0;
			32'd1506:
				output_byte = 8'd0;
			32'd1507:
				output_byte = 8'd4;
			32'd1508:
				output_byte = 8'd1;
			32'd1509:
				output_byte = 8'd0;
			32'd1510:
				output_byte = 8'd0;
			32'd1511:
				output_byte = 8'd0;
			32'd1512:
				output_byte = 8'd2;
			32'd1513:
				output_byte = 8'd0;
			32'd1514:
				output_byte = 8'd0;
			32'd1515:
				output_byte = 8'd0;
			32'd1516:
				output_byte = 8'd2;
			32'd1517:
				output_byte = 8'd1;
			32'd1518:
				output_byte = 8'd0;
			32'd1519:
				output_byte = 8'd0;
			32'd1520:
				output_byte = 8'd0;
			32'd1521:
				output_byte = 8'd0;
			32'd1522:
				output_byte = 8'd0;
			32'd1523:
				output_byte = 8'd0;
			32'd1524:
				output_byte = 8'd0;
			32'd1525:
				output_byte = 8'd20;
			32'd1526:
				output_byte = 8'd0;
			32'd1527:
				output_byte = 8'd0;
			32'd1528:
				output_byte = 8'd0;
			32'd1529:
				output_byte = 8'd0;
			32'd1530:
				output_byte = 8'd1;
			32'd1531:
				output_byte = 8'd0;
			32'd1532:
				output_byte = 8'd0;
			32'd1533:
				output_byte = 8'd0;
			32'd1534:
				output_byte = 8'd1;
			32'd1535:
				output_byte = 8'd44;
			32'd1536:
				output_byte = 8'd0;
			32'd1537:
				output_byte = 8'd0;
			32'd1538:
				output_byte = 8'd0;
			32'd1539:
				output_byte = 8'd2;
			32'd1540:
				output_byte = 8'd0;
			32'd1541:
				output_byte = 8'd0;
			32'd1542:
				output_byte = 8'd0;
			32'd1543:
				output_byte = 8'd3;
			32'd1544:
				output_byte = 8'd1;
			32'd1545:
				output_byte = 8'd0;
			32'd1546:
				output_byte = 8'd0;
			32'd1547:
				output_byte = 8'd0;
			32'd1548:
				output_byte = 8'd2;
			32'd1549:
				output_byte = 8'd0;
			32'd1550:
				output_byte = 8'd0;
			32'd1551:
				output_byte = 8'd0;
			32'd1552:
				output_byte = 8'd20;
			32'd1553:
				output_byte = 8'd48;
			32'd1554:
				output_byte = 8'd0;
			32'd1555:
				output_byte = 8'd0;
			32'd1556:
				output_byte = 8'd0;
			32'd1557:
				output_byte = 8'd2;
			32'd1558:
				output_byte = 8'd0;
			32'd1559:
				output_byte = 8'd0;
			32'd1560:
				output_byte = 8'd0;
			32'd1561:
				output_byte = 8'd3;
			32'd1562:
				output_byte = 8'd1;
			32'd1563:
				output_byte = 8'd0;
			32'd1564:
				output_byte = 8'd0;
			32'd1565:
				output_byte = 8'd0;
			32'd1566:
				output_byte = 8'd2;
			32'd1567:
				output_byte = 8'd0;
			32'd1568:
				output_byte = 8'd0;
			32'd1569:
				output_byte = 8'd0;
			32'd1570:
				output_byte = 8'd2;
			32'd1571:
				output_byte = 8'd1;
			32'd1572:
				output_byte = 8'd0;
			32'd1573:
				output_byte = 8'd0;
			32'd1574:
				output_byte = 8'd0;
			32'd1575:
				output_byte = 8'd4;
			32'd1576:
				output_byte = 8'd0;
			32'd1577:
				output_byte = 8'd0;
			32'd1578:
				output_byte = 8'd0;
			32'd1579:
				output_byte = 8'd1;
			32'd1580:
				output_byte = 8'd0;
			32'd1581:
				output_byte = 8'd0;
			32'd1582:
				output_byte = 8'd0;
			32'd1583:
				output_byte = 8'd0;
			32'd1584:
				output_byte = 8'd1;
			32'd1585:
				output_byte = 8'd0;
			32'd1586:
				output_byte = 8'd0;
			32'd1587:
				output_byte = 8'd0;
			32'd1588:
				output_byte = 8'd1;
			32'd1589:
				output_byte = 8'd4;
			32'd1590:
				output_byte = 8'd0;
			32'd1591:
				output_byte = 8'd0;
			32'd1592:
				output_byte = 8'd0;
			32'd1593:
				output_byte = 8'd2;
			32'd1594:
				output_byte = 8'd0;
			32'd1595:
				output_byte = 8'd0;
			32'd1596:
				output_byte = 8'd0;
			32'd1597:
				output_byte = 8'd5;
			32'd1598:
				output_byte = 8'd1;
			32'd1599:
				output_byte = 8'd0;
			32'd1600:
				output_byte = 8'd0;
			32'd1601:
				output_byte = 8'd0;
			32'd1602:
				output_byte = 8'd2;
			32'd1603:
				output_byte = 8'd0;
			32'd1604:
				output_byte = 8'd0;
			32'd1605:
				output_byte = 8'd0;
			32'd1606:
				output_byte = 8'd20;
			32'd1607:
				output_byte = 8'd0;
			32'd1608:
				output_byte = 8'd0;
			32'd1609:
				output_byte = 8'd0;
			32'd1610:
				output_byte = 8'd0;
			32'd1611:
				output_byte = 8'd1;
			32'd1612:
				output_byte = 8'd0;
			32'd1613:
				output_byte = 8'd0;
			32'd1614:
				output_byte = 8'd0;
			32'd1615:
				output_byte = 8'd1;
			32'd1616:
				output_byte = 8'd36;
			32'd1617:
				output_byte = 8'd0;
			32'd1618:
				output_byte = 8'd0;
			32'd1619:
				output_byte = 8'd0;
			32'd1620:
				output_byte = 8'd2;
			32'd1621:
				output_byte = 8'd0;
			32'd1622:
				output_byte = 8'd0;
			32'd1623:
				output_byte = 8'd0;
			32'd1624:
				output_byte = 8'd3;
			32'd1625:
				output_byte = 8'd1;
			32'd1626:
				output_byte = 8'd0;
			32'd1627:
				output_byte = 8'd0;
			32'd1628:
				output_byte = 8'd0;
			32'd1629:
				output_byte = 8'd2;
			32'd1630:
				output_byte = 8'd0;
			32'd1631:
				output_byte = 8'd0;
			32'd1632:
				output_byte = 8'd0;
			32'd1633:
				output_byte = 8'd20;
			32'd1634:
				output_byte = 8'd1;
			32'd1635:
				output_byte = 8'd0;
			32'd1636:
				output_byte = 8'd0;
			32'd1637:
				output_byte = 8'd0;
			32'd1638:
				output_byte = 8'd2;
			32'd1639:
				output_byte = 8'd0;
			32'd1640:
				output_byte = 8'd0;
			32'd1641:
				output_byte = 8'd0;
			32'd1642:
				output_byte = 8'd4;
			32'd1643:
				output_byte = 8'd1;
			32'd1644:
				output_byte = 8'd0;
			32'd1645:
				output_byte = 8'd0;
			32'd1646:
				output_byte = 8'd0;
			32'd1647:
				output_byte = 8'd2;
			32'd1648:
				output_byte = 8'd0;
			32'd1649:
				output_byte = 8'd0;
			32'd1650:
				output_byte = 8'd0;
			32'd1651:
				output_byte = 8'd2;
			32'd1652:
				output_byte = 8'd1;
			32'd1653:
				output_byte = 8'd0;
			32'd1654:
				output_byte = 8'd0;
			32'd1655:
				output_byte = 8'd0;
			32'd1656:
				output_byte = 8'd36;
			32'd1657:
				output_byte = 8'd0;
			32'd1658:
				output_byte = 8'd0;
			32'd1659:
				output_byte = 8'd0;
			32'd1660:
				output_byte = 8'd20;
			32'd1661:
				output_byte = 8'd0;
			32'd1662:
				output_byte = 8'd0;
			32'd1663:
				output_byte = 8'd0;
			32'd1664:
				output_byte = 8'd0;
			32'd1665:
				output_byte = 8'd1;
			32'd1666:
				output_byte = 8'd0;
			32'd1667:
				output_byte = 8'd0;
			32'd1668:
				output_byte = 8'd0;
			32'd1669:
				output_byte = 8'd1;
			32'd1670:
				output_byte = 8'd40;
			32'd1671:
				output_byte = 8'd0;
			32'd1672:
				output_byte = 8'd0;
			32'd1673:
				output_byte = 8'd0;
			32'd1674:
				output_byte = 8'd2;
			32'd1675:
				output_byte = 8'd0;
			32'd1676:
				output_byte = 8'd0;
			32'd1677:
				output_byte = 8'd0;
			32'd1678:
				output_byte = 8'd3;
			32'd1679:
				output_byte = 8'd1;
			32'd1680:
				output_byte = 8'd0;
			32'd1681:
				output_byte = 8'd0;
			32'd1682:
				output_byte = 8'd0;
			32'd1683:
				output_byte = 8'd2;
			32'd1684:
				output_byte = 8'd0;
			32'd1685:
				output_byte = 8'd0;
			32'd1686:
				output_byte = 8'd0;
			32'd1687:
				output_byte = 8'd20;
			32'd1688:
				output_byte = 8'd10;
			32'd1689:
				output_byte = 8'd0;
			32'd1690:
				output_byte = 8'd0;
			32'd1691:
				output_byte = 8'd0;
			32'd1692:
				output_byte = 8'd2;
			32'd1693:
				output_byte = 8'd0;
			32'd1694:
				output_byte = 8'd0;
			32'd1695:
				output_byte = 8'd0;
			32'd1696:
				output_byte = 8'd22;
			32'd1697:
				output_byte = 8'd1;
			32'd1698:
				output_byte = 8'd0;
			32'd1699:
				output_byte = 8'd0;
			32'd1700:
				output_byte = 8'd0;
			32'd1701:
				output_byte = 8'd2;
			32'd1702:
				output_byte = 8'd0;
			32'd1703:
				output_byte = 8'd0;
			32'd1704:
				output_byte = 8'd0;
			32'd1705:
				output_byte = 8'd2;
			32'd1706:
				output_byte = 8'd1;
			32'd1707:
				output_byte = 8'd0;
			32'd1708:
				output_byte = 8'd0;
			32'd1709:
				output_byte = 8'd0;
			32'd1710:
				output_byte = 8'd40;
			32'd1711:
				output_byte = 8'd0;
			32'd1712:
				output_byte = 8'd0;
			32'd1713:
				output_byte = 8'd0;
			32'd1714:
				output_byte = 8'd8;
			32'd1715:
				output_byte = 8'd1;
			32'd1716:
				output_byte = 8'd0;
			32'd1717:
				output_byte = 8'd0;
			32'd1718:
				output_byte = 8'd0;
			32'd1719:
				output_byte = 8'd1;
			32'd1720:
				output_byte = 8'd0;
			32'd1721:
				output_byte = 8'd0;
			32'd1722:
				output_byte = 8'd0;
			32'd1723:
				output_byte = 8'd10;
			32'd1724:
				output_byte = 8'd155;
			32'd1725:
				output_byte = 8'd4;
			32'd1726:
				output_byte = 8'd0;
			32'd1727:
				output_byte = 8'd0;
			32'd1728:
				output_byte = 8'd0;
			32'd1729:
				output_byte = 8'd0;
			32'd1730:
				output_byte = 8'd0;
			32'd1731:
				output_byte = 8'd0;
			32'd1732:
				output_byte = 8'd20;
			32'd1733:
				output_byte = 8'd0;
			32'd1734:
				output_byte = 8'd0;
			32'd1735:
				output_byte = 8'd0;
			32'd1736:
				output_byte = 8'd0;
			32'd1737:
				output_byte = 8'd1;
			32'd1738:
				output_byte = 8'd0;
			32'd1739:
				output_byte = 8'd0;
			32'd1740:
				output_byte = 8'd0;
			32'd1741:
				output_byte = 8'd1;
			32'd1742:
				output_byte = 8'd12;
			32'd1743:
				output_byte = 8'd0;
			32'd1744:
				output_byte = 8'd0;
			32'd1745:
				output_byte = 8'd0;
			32'd1746:
				output_byte = 8'd2;
			32'd1747:
				output_byte = 8'd0;
			32'd1748:
				output_byte = 8'd0;
			32'd1749:
				output_byte = 8'd0;
			32'd1750:
				output_byte = 8'd3;
			32'd1751:
				output_byte = 8'd1;
			32'd1752:
				output_byte = 8'd0;
			32'd1753:
				output_byte = 8'd0;
			32'd1754:
				output_byte = 8'd0;
			32'd1755:
				output_byte = 8'd2;
			32'd1756:
				output_byte = 8'd0;
			32'd1757:
				output_byte = 8'd0;
			32'd1758:
				output_byte = 8'd0;
			32'd1759:
				output_byte = 8'd20;
			32'd1760:
				output_byte = 8'd1;
			32'd1761:
				output_byte = 8'd0;
			32'd1762:
				output_byte = 8'd0;
			32'd1763:
				output_byte = 8'd0;
			32'd1764:
				output_byte = 8'd2;
			32'd1765:
				output_byte = 8'd0;
			32'd1766:
				output_byte = 8'd0;
			32'd1767:
				output_byte = 8'd0;
			32'd1768:
				output_byte = 8'd3;
			32'd1769:
				output_byte = 8'd1;
			32'd1770:
				output_byte = 8'd0;
			32'd1771:
				output_byte = 8'd0;
			32'd1772:
				output_byte = 8'd0;
			32'd1773:
				output_byte = 8'd2;
			32'd1774:
				output_byte = 8'd0;
			32'd1775:
				output_byte = 8'd0;
			32'd1776:
				output_byte = 8'd0;
			32'd1777:
				output_byte = 8'd2;
			32'd1778:
				output_byte = 8'd1;
			32'd1779:
				output_byte = 8'd0;
			32'd1780:
				output_byte = 8'd0;
			32'd1781:
				output_byte = 8'd0;
			32'd1782:
				output_byte = 8'd12;
			32'd1783:
				output_byte = 8'd0;
			32'd1784:
				output_byte = 8'd0;
			32'd1785:
				output_byte = 8'd0;
			32'd1786:
				output_byte = 8'd20;
			32'd1787:
				output_byte = 8'd0;
			32'd1788:
				output_byte = 8'd0;
			32'd1789:
				output_byte = 8'd0;
			32'd1790:
				output_byte = 8'd0;
			32'd1791:
				output_byte = 8'd1;
			32'd1792:
				output_byte = 8'd0;
			32'd1793:
				output_byte = 8'd0;
			32'd1794:
				output_byte = 8'd0;
			32'd1795:
				output_byte = 8'd1;
			32'd1796:
				output_byte = 8'd16;
			32'd1797:
				output_byte = 8'd0;
			32'd1798:
				output_byte = 8'd0;
			32'd1799:
				output_byte = 8'd0;
			32'd1800:
				output_byte = 8'd2;
			32'd1801:
				output_byte = 8'd0;
			32'd1802:
				output_byte = 8'd0;
			32'd1803:
				output_byte = 8'd0;
			32'd1804:
				output_byte = 8'd3;
			32'd1805:
				output_byte = 8'd1;
			32'd1806:
				output_byte = 8'd0;
			32'd1807:
				output_byte = 8'd0;
			32'd1808:
				output_byte = 8'd0;
			32'd1809:
				output_byte = 8'd2;
			32'd1810:
				output_byte = 8'd0;
			32'd1811:
				output_byte = 8'd0;
			32'd1812:
				output_byte = 8'd0;
			32'd1813:
				output_byte = 8'd20;
			32'd1814:
				output_byte = 8'd1;
			32'd1815:
				output_byte = 8'd0;
			32'd1816:
				output_byte = 8'd0;
			32'd1817:
				output_byte = 8'd0;
			32'd1818:
				output_byte = 8'd2;
			32'd1819:
				output_byte = 8'd0;
			32'd1820:
				output_byte = 8'd0;
			32'd1821:
				output_byte = 8'd0;
			32'd1822:
				output_byte = 8'd3;
			32'd1823:
				output_byte = 8'd1;
			32'd1824:
				output_byte = 8'd0;
			32'd1825:
				output_byte = 8'd0;
			32'd1826:
				output_byte = 8'd0;
			32'd1827:
				output_byte = 8'd2;
			32'd1828:
				output_byte = 8'd0;
			32'd1829:
				output_byte = 8'd0;
			32'd1830:
				output_byte = 8'd0;
			32'd1831:
				output_byte = 8'd2;
			32'd1832:
				output_byte = 8'd1;
			32'd1833:
				output_byte = 8'd0;
			32'd1834:
				output_byte = 8'd0;
			32'd1835:
				output_byte = 8'd0;
			32'd1836:
				output_byte = 8'd16;
			32'd1837:
				output_byte = 8'd0;
			32'd1838:
				output_byte = 8'd0;
			32'd1839:
				output_byte = 8'd0;
			32'd1840:
				output_byte = 8'd8;
			32'd1841:
				output_byte = 8'd1;
			32'd1842:
				output_byte = 8'd0;
			32'd1843:
				output_byte = 8'd0;
			32'd1844:
				output_byte = 8'd0;
			32'd1845:
				output_byte = 8'd1;
			32'd1846:
				output_byte = 8'd0;
			32'd1847:
				output_byte = 8'd0;
			32'd1848:
				output_byte = 8'd0;
			32'd1849:
				output_byte = 8'd10;
			32'd1850:
				output_byte = 8'd126;
			32'd1851:
				output_byte = 8'd0;
			32'd1852:
				output_byte = 8'd0;
			32'd1853:
				output_byte = 8'd0;
			32'd1854:
				output_byte = 8'd0;
			32'd1855:
				output_byte = 8'd0;
			32'd1856:
				output_byte = 8'd0;
			32'd1857:
				output_byte = 8'd0;
			32'd1858:
				output_byte = 8'd13;
			32'd1859:
				output_byte = 8'd0;
			32'd1860:
				output_byte = 8'd0;
			32'd1861:
				output_byte = 8'd0;
			32'd1862:
				output_byte = 8'd0;
			32'd1863:
				output_byte = 8'd0;
			32'd1864:
				output_byte = 8'd0;
			32'd1865:
				output_byte = 8'd0;
			32'd1866:
				output_byte = 8'd0;
			default:
				output_byte = 8'd0;
		endcase
	end
endmodule