module rom(input[31:0] address, output reg [7:0] output_byte, output done);
	assign done = (address == 32'd231) ? 1'b1 : 1'b0;
	always @(address)
	begin
		case (address)
			32'd0:
				output_byte = 8'd1;
			32'd1:
				output_byte = 8'd0;
			32'd2:
				output_byte = 8'd0;
			32'd3:
				output_byte = 8'd0;
			32'd4:
				output_byte = 8'd1;
			32'd5:
				output_byte = 8'd0;
			32'd6:
				output_byte = 8'd0;
			32'd7:
				output_byte = 8'd0;
			32'd8:
				output_byte = 8'd0;
			32'd9:
				output_byte = 8'd0;
			32'd10:
				output_byte = 8'd0;
			32'd11:
				output_byte = 8'd0;
			32'd12:
				output_byte = 8'd1;
			32'd13:
				output_byte = 8'd0;
			32'd14:
				output_byte = 8'd0;
			32'd15:
				output_byte = 8'd0;
			32'd16:
				output_byte = 8'd17;
			32'd17:
				output_byte = 8'd0;
			32'd18:
				output_byte = 8'd0;
			32'd19:
				output_byte = 8'd0;
			32'd20:
				output_byte = 8'd32;
			32'd21:
				output_byte = 8'd161;
			32'd22:
				output_byte = 8'd7;
			32'd23:
				output_byte = 8'd0;
			32'd24:
				output_byte = 8'd14;
			32'd25:
				output_byte = 8'd1;
			32'd26:
				output_byte = 8'd0;
			32'd27:
				output_byte = 8'd0;
			32'd28:
				output_byte = 8'd0;
			32'd29:
				output_byte = 8'd0;
			32'd30:
				output_byte = 8'd2;
			32'd31:
				output_byte = 8'd0;
			32'd32:
				output_byte = 8'd0;
			32'd33:
				output_byte = 8'd0;
			32'd34:
				output_byte = 8'd1;
			32'd35:
				output_byte = 8'd4;
			32'd36:
				output_byte = 8'd0;
			32'd37:
				output_byte = 8'd0;
			32'd38:
				output_byte = 8'd0;
			32'd39:
				output_byte = 8'd3;
			32'd40:
				output_byte = 8'd0;
			32'd41:
				output_byte = 8'd0;
			32'd42:
				output_byte = 8'd0;
			32'd43:
				output_byte = 8'd1;
			32'd44:
				output_byte = 8'd8;
			32'd45:
				output_byte = 8'd0;
			32'd46:
				output_byte = 8'd0;
			32'd47:
				output_byte = 8'd0;
			32'd48:
				output_byte = 8'd4;
			32'd49:
				output_byte = 8'd0;
			32'd50:
				output_byte = 8'd0;
			32'd51:
				output_byte = 8'd0;
			32'd52:
				output_byte = 8'd1;
			32'd53:
				output_byte = 8'd16;
			32'd54:
				output_byte = 8'd0;
			32'd55:
				output_byte = 8'd0;
			32'd56:
				output_byte = 8'd0;
			32'd57:
				output_byte = 8'd5;
			32'd58:
				output_byte = 8'd0;
			32'd59:
				output_byte = 8'd0;
			32'd60:
				output_byte = 8'd0;
			32'd61:
				output_byte = 8'd1;
			32'd62:
				output_byte = 8'd12;
			32'd63:
				output_byte = 8'd0;
			32'd64:
				output_byte = 8'd0;
			32'd65:
				output_byte = 8'd0;
			32'd66:
				output_byte = 8'd6;
			32'd67:
				output_byte = 8'd0;
			32'd68:
				output_byte = 8'd0;
			32'd69:
				output_byte = 8'd0;
			32'd70:
				output_byte = 8'd1;
			32'd71:
				output_byte = 8'd20;
			32'd72:
				output_byte = 8'd0;
			32'd73:
				output_byte = 8'd0;
			32'd74:
				output_byte = 8'd0;
			32'd75:
				output_byte = 8'd7;
			32'd76:
				output_byte = 8'd0;
			32'd77:
				output_byte = 8'd0;
			32'd78:
				output_byte = 8'd0;
			32'd79:
				output_byte = 8'd4;
			32'd80:
				output_byte = 8'd7;
			32'd81:
				output_byte = 8'd0;
			32'd82:
				output_byte = 8'd0;
			32'd83:
				output_byte = 8'd0;
			32'd84:
				output_byte = 8'd6;
			32'd85:
				output_byte = 8'd0;
			32'd86:
				output_byte = 8'd0;
			32'd87:
				output_byte = 8'd0;
			32'd88:
				output_byte = 8'd7;
			32'd89:
				output_byte = 8'd1;
			32'd90:
				output_byte = 8'd0;
			32'd91:
				output_byte = 8'd0;
			32'd92:
				output_byte = 8'd0;
			32'd93:
				output_byte = 8'd7;
			32'd94:
				output_byte = 8'd0;
			32'd95:
				output_byte = 8'd0;
			32'd96:
				output_byte = 8'd0;
			32'd97:
				output_byte = 8'd8;
			32'd98:
				output_byte = 8'd7;
			32'd99:
				output_byte = 8'd0;
			32'd100:
				output_byte = 8'd0;
			32'd101:
				output_byte = 8'd0;
			32'd102:
				output_byte = 8'd6;
			32'd103:
				output_byte = 8'd0;
			32'd104:
				output_byte = 8'd0;
			32'd105:
				output_byte = 8'd0;
			32'd106:
				output_byte = 8'd10;
			32'd107:
				output_byte = 8'd99;
			32'd108:
				output_byte = 8'd0;
			32'd109:
				output_byte = 8'd0;
			32'd110:
				output_byte = 8'd0;
			32'd111:
				output_byte = 8'd0;
			32'd112:
				output_byte = 8'd0;
			32'd113:
				output_byte = 8'd0;
			32'd114:
				output_byte = 8'd0;
			32'd115:
				output_byte = 8'd11;
			32'd116:
				output_byte = 8'd54;
			32'd117:
				output_byte = 8'd0;
			32'd118:
				output_byte = 8'd0;
			32'd119:
				output_byte = 8'd0;
			32'd120:
				output_byte = 8'd0;
			32'd121:
				output_byte = 8'd0;
			32'd122:
				output_byte = 8'd0;
			32'd123:
				output_byte = 8'd0;
			32'd124:
				output_byte = 8'd1;
			32'd125:
				output_byte = 8'd20;
			32'd126:
				output_byte = 8'd0;
			32'd127:
				output_byte = 8'd0;
			32'd128:
				output_byte = 8'd0;
			32'd129:
				output_byte = 8'd7;
			32'd130:
				output_byte = 8'd0;
			32'd131:
				output_byte = 8'd0;
			32'd132:
				output_byte = 8'd0;
			32'd133:
				output_byte = 8'd3;
			32'd134:
				output_byte = 8'd2;
			32'd135:
				output_byte = 8'd0;
			32'd136:
				output_byte = 8'd0;
			32'd137:
				output_byte = 8'd0;
			32'd138:
				output_byte = 8'd3;
			32'd139:
				output_byte = 8'd0;
			32'd140:
				output_byte = 8'd0;
			32'd141:
				output_byte = 8'd0;
			32'd142:
				output_byte = 8'd7;
			32'd143:
				output_byte = 8'd3;
			32'd144:
				output_byte = 8'd0;
			32'd145:
				output_byte = 8'd0;
			32'd146:
				output_byte = 8'd0;
			32'd147:
				output_byte = 8'd2;
			32'd148:
				output_byte = 8'd0;
			32'd149:
				output_byte = 8'd0;
			32'd150:
				output_byte = 8'd0;
			32'd151:
				output_byte = 8'd7;
			32'd152:
				output_byte = 8'd1;
			32'd153:
				output_byte = 8'd0;
			32'd154:
				output_byte = 8'd0;
			32'd155:
				output_byte = 8'd0;
			32'd156:
				output_byte = 8'd3;
			32'd157:
				output_byte = 8'd0;
			32'd158:
				output_byte = 8'd0;
			32'd159:
				output_byte = 8'd0;
			32'd160:
				output_byte = 8'd5;
			32'd161:
				output_byte = 8'd3;
			32'd162:
				output_byte = 8'd0;
			32'd163:
				output_byte = 8'd0;
			32'd164:
				output_byte = 8'd0;
			32'd165:
				output_byte = 8'd0;
			32'd166:
				output_byte = 8'd0;
			32'd167:
				output_byte = 8'd0;
			32'd168:
				output_byte = 8'd0;
			32'd169:
				output_byte = 8'd3;
			32'd170:
				output_byte = 8'd4;
			32'd171:
				output_byte = 8'd0;
			32'd172:
				output_byte = 8'd0;
			32'd173:
				output_byte = 8'd0;
			32'd174:
				output_byte = 8'd6;
			32'd175:
				output_byte = 8'd0;
			32'd176:
				output_byte = 8'd0;
			32'd177:
				output_byte = 8'd0;
			32'd178:
				output_byte = 8'd7;
			32'd179:
				output_byte = 8'd1;
			32'd180:
				output_byte = 8'd0;
			32'd181:
				output_byte = 8'd0;
			32'd182:
				output_byte = 8'd0;
			32'd183:
				output_byte = 8'd4;
			32'd184:
				output_byte = 8'd0;
			32'd185:
				output_byte = 8'd0;
			32'd186:
				output_byte = 8'd0;
			32'd187:
				output_byte = 8'd8;
			32'd188:
				output_byte = 8'd4;
			32'd189:
				output_byte = 8'd0;
			32'd190:
				output_byte = 8'd0;
			32'd191:
				output_byte = 8'd0;
			32'd192:
				output_byte = 8'd5;
			32'd193:
				output_byte = 8'd0;
			32'd194:
				output_byte = 8'd0;
			32'd195:
				output_byte = 8'd0;
			32'd196:
				output_byte = 8'd9;
			32'd197:
				output_byte = 8'd54;
			32'd198:
				output_byte = 8'd0;
			32'd199:
				output_byte = 8'd0;
			32'd200:
				output_byte = 8'd0;
			32'd201:
				output_byte = 8'd0;
			32'd202:
				output_byte = 8'd0;
			32'd203:
				output_byte = 8'd0;
			32'd204:
				output_byte = 8'd0;
			32'd205:
				output_byte = 8'd10;
			32'd206:
				output_byte = 8'd54;
			32'd207:
				output_byte = 8'd0;
			32'd208:
				output_byte = 8'd0;
			32'd209:
				output_byte = 8'd0;
			32'd210:
				output_byte = 8'd0;
			32'd211:
				output_byte = 8'd0;
			32'd212:
				output_byte = 8'd0;
			32'd213:
				output_byte = 8'd0;
			32'd214:
				output_byte = 8'd11;
			32'd215:
				output_byte = 8'd198;
			32'd216:
				output_byte = 8'd0;
			32'd217:
				output_byte = 8'd0;
			32'd218:
				output_byte = 8'd0;
			32'd219:
				output_byte = 8'd0;
			32'd220:
				output_byte = 8'd0;
			32'd221:
				output_byte = 8'd0;
			32'd222:
				output_byte = 8'd0;
			32'd223:
				output_byte = 8'd13;
			32'd224:
				output_byte = 8'd0;
			32'd225:
				output_byte = 8'd0;
			32'd226:
				output_byte = 8'd0;
			32'd227:
				output_byte = 8'd0;
			32'd228:
				output_byte = 8'd0;
			32'd229:
				output_byte = 8'd0;
			32'd230:
				output_byte = 8'd0;
			32'd231:
				output_byte = 8'd0;
			default:
				output_byte = 8'd0;
		endcase
	end
endmodule